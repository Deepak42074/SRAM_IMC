* NGSPICE file created from Integrated_bitcell_with_dummy_cells_flat.ext - technology: sky130B

.subckt Integrated_bitcell_with_dummy_cells_flat PRE_SRAM RWL[0] WWL[0] RWLB[0] RWL[1]
+ WWL[1] RWLB[1] RWL[2] WWL[2] RWLB[2] RWL[3] WWL[3] RWLB[3] RWL[4] WWL[4] RWLB[4]
+ RWL[5] WWL[5] RWLB[5] RWL[6] WWL[6] RWLB[6] RWL[7] WWL[7] RWLB[7] RWL[8] WWL[8]
+ RWLB[8] RWL[9] WWL[9] RWLB[9] RWL[10] WWL[10] RWLB[10] RWL[11] WWL[11] RWLB[11]
+ RWL[12] WWL[12] RWLB[12] RWL[13] WWL[13] RWLB[13] RWL[14] WWL[14] RWLB[14] RWL[15]
+ WWL[15] RWLB[15] PRE_VLSA WE PRE_CLSA VCLP SAEN ADC0_OUT[0] ADC0_OUT[1] ADC0_OUT[2]
+ ADC0_OUT[3] ADC1_OUT[0] ADC1_OUT[1] ADC1_OUT[2] ADC1_OUT[3] ADC2_OUT[0] ADC2_OUT[1]
+ ADC2_OUT[2] ADC2_OUT[3] ADC3_OUT[0] ADC3_OUT[1] ADC3_OUT[2] ADC3_OUT[3] ADC4_OUT[0]
+ ADC4_OUT[1] ADC4_OUT[2] ADC4_OUT[3] ADC5_OUT[0] ADC5_OUT[1] ADC5_OUT[2] ADC5_OUT[3]
+ ADC6_OUT[0] ADC6_OUT[1] ADC6_OUT[2] ADC6_OUT[3] ADC7_OUT[0] ADC7_OUT[1] ADC7_OUT[2]
+ ADC7_OUT[3] ADC8_OUT[0] ADC8_OUT[1] ADC8_OUT[2] ADC8_OUT[3] ADC9_OUT[0] ADC9_OUT[1]
+ ADC9_OUT[2] ADC9_OUT[3] ADC10_OUT[0] ADC10_OUT[1] ADC10_OUT[2] ADC10_OUT[3] ADC11_OUT[0]
+ ADC11_OUT[1] ADC11_OUT[2] ADC11_OUT[3] ADC12_OUT[0] ADC12_OUT[1] ADC12_OUT[2] ADC12_OUT[3]
+ ADC13_OUT[0] ADC13_OUT[1] ADC13_OUT[2] ADC13_OUT[3] ADC14_OUT[0] ADC14_OUT[1] ADC14_OUT[2]
+ ADC14_OUT[3] ADC15_OUT[0] ADC15_OUT[1] ADC15_OUT[2] ADC15_OUT[3] Din[0] Din[1] Din[2]
+ Din[3] Din[4] Din[5] Din[6] Din[7] Din[8] Din[9] Din[10] Din[11] Din[12] Din[13]
+ Din[14] Din[15] WWLD[0] WWLD[1] WWLD[2] WWLD[3] WWLD[4] WWLD[5] WWLD[6] WWLD[7]
+ SA_OUT[0] SA_OUT[1] SA_OUT[2] SA_OUT[3] SA_OUT[4] SA_OUT[5] SA_OUT[6] SA_OUT[7]
+ SA_OUT[8] SA_OUT[9] SA_OUT[10] SA_OUT[11] SA_OUT[12] SA_OUT[13] SA_OUT[14] SA_OUT[15]
+ EN PRE_A Iref0 Iref1 Iref2 Iref3 VSS VDD
X0 a_2015_2180.t0 a_2002_2165.t3 VSS.t1274 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 SA_OUT[5].t0 PRE_VLSA.t0 VDD.t1167 VDD.t1166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 a_8340_n953.t11 VSS.t764 a_8340_n812.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VSS.t397 a_3247_3666.t3 a_3617_3666.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VSS.t389 a_4397_1698.t3 a_4767_1698.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_1440_452.t0 a_1427_437.t3 VSS.t393 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_372_1216.t1 a_277_1201.t3 VSS.t253 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VSS.t403 a_7827_n2234.t2 a_7950_n2132.t0 VSS.t402 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VSS.t391 a_3247_n512.t3 a_3152_n527.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_2097_4148.t1 a_2002_4133.t3 VDD.t311 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_8422_3184.t1 a_8327_3169.t3 VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_3247_2180.t1 a_3152_2165.t3 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VDD.t1165 PRE_VLSA.t1 a_2035_n1371.t2 VDD.t1164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X13 a_865_n953.t6 VSS.t763 a_865_n812.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_3740_n953.t9 VSS.t762 a_3740_4686.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_8792_3425.t1 RWLB[1].t0 a_8340_n953.t2 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VSS.t228 a_4972_1698.t3 a_4877_1683.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_8422_n30.t0 a_8327_n45.t3 VSS.t244 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X18 a_8221_n7216.t1 ADC10_OUT[2].t3 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 VSS.t158 a_4397_n812.t3 a_4767_n812.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_2577_3410.t0 WWL[1].t0 a_2845_4887.t3 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_3822_693.t1 a_3727_678.t3 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VSS.t263 SAEN.t0 a_n3792_n8026.t1 VSS.t262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X23 a_n52_n8583.t0 PRE_CLSA.t0 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 VSS.t108 a_4972_n812.t3 a_4877_n827.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_3042_4445.t0 VSS.t761 a_2590_n953.t4 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_5547_211.t1 a_5452_196.t3 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VDD.t65 a_2672_n30.t3 a_2577_n45.t1 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VSS.t104 a_6697_n271.t3 a_6602_n286.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_4315_n953.t5 VSS.t760 a_4315_4445.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 SA_OUT[10].t2 PRE_VLSA.t2 VDD.t1163 VDD.t1162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X31 a_7190_n953.t7 VSS.t759 a_7190_n512.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_4302_1201.t0 WWL[10].t0 a_4570_4887.t6 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_6615_975.t1 a_6602_960.t3 VSS.t112 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VSS.t3 a_n3827_n4378.t4 a_n3827_n7825.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X35 a_9613_n4470.t0 VCLP.t0 a_9475_n4470.t1 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X36 a_2084_n8026.t1 VCLP.t1 a_2049_n7825.t0 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X37 VSS.t100 a_4393_n2422.t4 a_4413_n7825.t1 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X38 VSS.t90 a_6697_3425.t3 a_6602_3410.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 a_8340_n953.t1 RWL[10].t0 a_8340_1216.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VSS.t84 a_947_452.t3 a_1317_452.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_5465_2662.t0 a_5452_2647.t3 VSS.t79 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 VDD.t89 PRE_CLSA.t1 ADC13_OUT[2].t2 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 a_7752_3892.t0 WWLD[3].t0 a_8020_4887.t5 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X44 a_290_n953.t26 RWL[0].t0 a_290_3666.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 a_6697_2180.t1 a_6602_2165.t3 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_865_n953.t2 RWL[10].t1 a_865_1216.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X47 VSS.t61 a_947_4445.t3 a_852_4430.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X48 VSS.t40 a_3822_3666.t3 a_4192_3666.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X49 VSS.t2416 a_4397_1216.t3 a_4767_1216.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 a_4877_1924.t0 WWL[7].t0 a_5145_4887.t5 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 a_1440_n512.t1 a_1427_n527.t3 VSS.t41 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X52 a_13864_n5850.t2 ADC15_OUT[1].t3 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X53 SA_OUT[7].t0 PRE_VLSA.t3 VDD.t1161 VDD.t1160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X54 VSS.t2363 a_3822_n512.t3 a_3727_n527.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X55 a_10797_n7203.t1 a_5743_n6391# a_10659_n7203.t2 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X56 VSS.t2402 a_8977_n2234.t2 a_9100_n2132.t0 VSS.t2401 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X57 VSS.t55 a_4972_1216.t3 a_4877_1201.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X58 VDD.t1159 PRE_VLSA.t4 a_3185_n1371.t0 VDD.t1158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 VSS.t2357 a_7847_3907.t3 a_8217_3907.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X60 VDD.t7 a_3822_975.t3 a_3727_960.t1 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X61 a_3247_2180.t0 a_3152_2165.t4 VSS.t109 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X62 VDD.t2185 a_4972_n1053.t3 a_4877_n1068.t1 VDD.t2184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X63 a_2015_n953.t23 RWL[2].t0 a_2015_3184.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X64 a_2590_n30.t1 a_2577_n45.t3 VSS.t110 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X65 a_4890_2421.t0 a_4877_2406.t3 VSS.t2173 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X66 a_7272_2421.t2 a_7177_2406.t3 VDD.t2176 VDD.t2175 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X67 a_6203_n2086.t0 WE.t0 a_6133_n953.t7 VSS.t2403 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 VSS.t2193 a_8997_n1053.t3 a_9367_n1053.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X69 a_3258_n953.t4 WWLD[3].t1 a_3247_3907.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X70 a_7177_3651.t0 WWL[0].t0 a_7445_4887.t14 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X71 a_4890_n271.t1 a_4877_n286.t3 VSS.t2353 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X72 a_7272_n271.t1 a_7177_n286.t3 VDD.t2160 VDD.t2159 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X73 VDD.t2154 a_2672_n512.t3 a_2577_n527.t2 VDD.t2153 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 VSS.t2188 a_8422_975.t3 a_8327_960.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X75 a_3247_n1053.t1 a_3152_n1068.t3 VDD.t1926 VDD.t1925 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 a_2672_n1053.t0 a_2577_n1068.t3 VSS.t2335 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X77 VDD.t329 a_3247_3666.t4 a_3152_3651.t2 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X78 a_8915_2662.t0 a_8902_2647.t3 VSS.t2343 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X79 VDD.t321 a_4397_1698.t4 a_4302_1683.t2 VDD.t320 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X80 SA_OUT[12].t0 PRE_VLSA.t5 VDD.t1157 VDD.t1156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X81 a_372_4445.t0 a_277_4430.t3 VSS.t2171 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X82 a_6040_2180.t0 a_6027_2165.t3 VSS.t2176 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X83 VSS.t2168 a_8422_1698.t3 a_8792_1698.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X84 a_7177_678.t0 WWL[12].t0 a_7445_4887.t16 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X85 a_3822_n812.t0 a_3727_n827.t3 VSS.t2161 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X86 VSS.t2333 a_7272_3666.t3 a_7642_3666.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X87 a_8327_1924.t0 WWL[7].t1 a_8595_4887.t7 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X88 VDD.t55 a_4397_n812.t4 a_4302_n827.t1 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X89 a_7752_3410.t0 WWL[1].t1 a_8020_4887.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X90 a_1440_n953.t18 RWL[3].t0 a_1440_2943.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 a_8902_1442.t0 WWL[9].t0 a_9170_4887.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X92 a_958_n953.t9 WWL[14].t0 a_947_211.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X93 VSS.t2250 a_7272_n512.t3 a_7177_n527.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X94 a_1317_4148.t0 VSS.t758 a_865_n953.t19 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X95 a_2672_2943.t2 a_2577_2928.t3 VDD.t1972 VDD.t1971 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X96 a_2467_2180.t0 RWLB[6].t0 a_2015_n953.t40 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 a_2683_n953.t17 WWL[0].t1 a_2672_3666.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 VSS.t2249 a_7847_n271.t3 a_8217_n271.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X99 VDD.t1978 a_7039_n8583.t3 ADC9_OUT[3].t2 VDD.t1977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X100 VSS.t265 SAEN.t1 a_3266_n3770.t0 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X101 a_9078_n2086.t0 WE.t1 a_9008_n953.t6 VSS.t2404 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 VSS.t2215 a_8422_n812.t3 a_8792_n812.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 VDD.t1960 a_4972_1457.t3 a_4877_1442.t2 VDD.t1959 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X104 a_3822_n30.t1 a_3727_n45.t3 VSS.t2218 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X105 a_n2207_n5338.t1 Iref1.t0 a_n2148_n5293.t1 VSS.t2219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X106 VSS.t2206 a_372_3666.t3 a_277_3651.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X107 VSS.t245 a_8422_n30.t3 a_8327_n45.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X108 a_1522_n1053.t1 a_1427_n1068.t3 VDD.t2130 VDD.t2129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 a_13171_n7203.t1 a_5743_n6391# a_13033_n7203.t1 VSS.t222 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X110 a_6697_2662.t0 a_6602_2647.t3 VSS.t2201 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X111 VSS.t2302 a_8997_1457.t3 a_9367_1457.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 a_3258_n953.t17 WWLD[4].t0 a_3247_n271.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 a_8997_n812.t1 a_8902_n827.t3 VDD.t2124 VDD.t2123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 a_4302_4430.t0 WWLD[1].t0 a_4570_4887.t15 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X115 VSS.t2204 a_7847_3425.t3 a_8217_3425.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 a_6708_n953.t4 WWLD[3].t2 a_6697_3907.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X117 a_6492_975.t0 RWLB[11].t0 a_6040_n953.t22 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X118 a_8340_n953.t21 VSS.t757 a_8340_4445.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X119 a_4408_n953.t1 WWL[11].t0 a_4397_975.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X120 a_545_4887.t8 WE.t2 a_593_n2086.t1 VSS.t2405 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 a_2672_n512.t1 a_2577_n527.t3 VSS.t2190 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X122 a_865_n953.t20 VSS.t756 a_865_4445.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X123 a_3258_n953.t0 WWL[1].t2 a_3247_3425.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X124 VSS.t2435 a_n1495_n4378.t4 a_n1495_n5092.t1 VSS.t2433 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X125 a_7858_n953.t14 WWLD[7].t0 a_7847_n1053.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X126 a_7765_452.t0 a_7752_437.t3 VSS.t2258 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 a_2519_n8071.t1 Iref3.t0 a_2578_n8026.t1 VSS.t1980 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X128 a_3493_n8583.t0 PRE_CLSA.t2 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X129 a_7353_n2086.t0 WE.t3 a_7283_n953.t7 VSS.t2406 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 VSS.t2454 a_2049_n4378.t0 a_2049_n4378.t1 VSS.t2453 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 VSS.t2428 a_4397_4445.t3 a_4767_4445.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X132 VDD.t2189 a_4397_1216.t4 a_4302_1201.t1 VDD.t2188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X133 a_3822_3907.t2 a_3727_3892.t3 VDD.t2211 VDD.t2210 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X134 a_947_452.t1 a_852_437.t3 VDD.t2209 VDD.t2208 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X135 a_4397_n1053.t1 a_4302_n1068.t3 VDD.t2219 VDD.t2218 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 a_3822_n1053.t1 a_3727_n1068.t3 VSS.t2311 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X137 VSS.t2441 a_4972_4445.t3 a_4877_4430.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X138 a_5917_2180.t0 RWLB[6].t1 a_5465_n953.t24 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X139 VDD.t2244 a_372_693.t3 a_277_678.t1 VDD.t2243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 VSS.t2483 a_8422_1216.t3 a_8792_1216.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X141 VDD.t2164 a_7847_3907.t4 a_7752_3892.t1 VDD.t2163 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 VDD.t2249 a_6122_452.t3 a_6027_437.t1 VDD.t2248 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X143 VSS.t2314 a_7843_n2422.t4 a_11514_n5092.t1 VSS.t2312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 VDD.t2245 a_9405_n7216.t3 ADC11_OUT[2].t2 VDD.t1655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 VDD.t2134 a_372_3907.t3 a_277_3892.t2 VDD.t2133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X146 a_2002_3169.t0 WWL[2].t0 a_2270_4887.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 a_6708_n953.t21 WWL[13].t0 a_6697_452.t1 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X148 a_372_n512.t2 a_277_n527.t3 VDD.t2000 VDD.t1999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X149 a_3740_n953.t45 RWL[4].t0 a_3740_2662.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X150 a_6708_n953.t7 WWLD[4].t1 a_6697_n271.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X151 VDD.t2156 a_8997_n1053.t4 a_8902_n1068.t1 VDD.t2155 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 a_3165_n953.t13 VSS.t755 a_3165_4148.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_6122_4148.t0 a_6027_4133.t3 VSS.t2480 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X154 a_6040_n953.t26 RWL[2].t1 a_6040_3184.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X155 a_7272_2180.t0 a_7177_2165.t3 VSS.t2472 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X156 a_2097_1698.t1 a_2002_1683.t3 VDD.t2234 VDD.t2233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X157 a_1892_n512.t0 VSS.t754 a_1440_n953.t17 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 VSS.t2257 a_8997_n30.t3 a_8902_n45.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X159 a_7283_n953.t5 WWLD[3].t3 a_7272_3907.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X160 a_7858_n953.t15 WWL[9].t1 a_7847_1457.t1 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 VSS.t1499 a_5632_n6430# a_13637_n6503.t1 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X162 a_6708_n953.t0 WWL[1].t3 a_6697_3425.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 a_3042_2421.t0 RWLB[5].t0 a_2590_n953.t47 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X164 a_6122_975.t2 a_6027_960.t3 VDD.t2004 VDD.t2003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X165 a_852_678.t0 WWL[12].t1 a_1120_4887.t7 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 a_6615_n953.t31 RWL[12].t0 a_6615_693.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X167 a_13864_n5850.t0 PRE_CLSA.t3 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X168 VDD.t2275 a_6697_n512.t3 a_6602_n527.t2 VDD.t2274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X169 VSS.t2525 a_2097_3184.t3 a_2467_3184.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X170 a_3042_n271.t0 VSS.t753 a_2590_n953.t3 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X171 a_3468_n2086.t1 a_3227_n2234.t2 VSS.t2505 VSS.t2504 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X172 VSS.t2487 a_5547_693.t3 a_5452_678.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X173 a_8902_4671.t0 WWLD[0].t0 a_9170_4887.t20 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X174 a_3165_3907.t1 a_3152_3892.t3 VSS.t2501 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X175 a_4315_n953.t48 RWL[5].t0 a_4315_2421.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X176 a_11549_n6503.t2 a_11776_n7216.t3 ADC13_OUT[2].t0 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X177 a_4448_n8026.t1 VCLP.t2 a_4413_n7825.t0 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X178 a_4397_693.t1 a_4302_678.t3 VSS.t2503 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X179 a_8340_n953.t48 RWL[14].t0 a_8340_211.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X180 a_5465_2943.t0 a_5452_2928.t3 VSS.t2292 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 a_7847_975.t2 a_7752_960.t3 VDD.t2255 VDD.t2254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X182 a_2577_678.t2 WWL[12].t2 a_2845_4887.t14 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X183 a_n3357_n7203.t0 VCLP.t3 a_n3495_n7203.t2 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X184 VDD.t1970 a_7847_n271.t4 a_7752_n286.t2 VDD.t1969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X185 a_10797_n4470.t0 VCLP.t4 a_10659_n4470.t1 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X186 VDD.t2257 a_4972_4686.t3 a_4877_4671.t1 VDD.t2256 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 a_3822_3425.t2 a_3727_3410.t3 VDD.t2265 VDD.t2264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X188 VSS.t153 a_7272_211.t3 a_7177_196.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X189 SA_OUT[2].t1 a_1460_n1371.t3 a_1703_n1770.t0 VSS.t154 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X190 a_6492_2180.t0 RWLB[6].t2 a_6040_n953.t23 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 VDD.t2010 a_372_n271.t3 a_277_n286.t1 VDD.t2009 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X192 a_11776_n4483.t1 ADC13_OUT[0].t3 VDD.t2106 VDD.t2105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X193 a_927_n2234.t1 Din[1].t0 VDD.t2287 VDD.t2286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X194 a_5342_4148.t0 VSS.t752 a_4890_n953.t16 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 a_n1233_n7216.t2 ADC2_OUT[2].t3 a_n1163_n7203.t2 VSS.t1879 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X196 VSS.t2289 a_8997_4686.t3 a_9367_4686.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X197 a_5452_3169.t2 WWL[2].t1 a_5720_4887.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X198 VDD.t2128 a_8997_1457.t4 a_8902_1442.t1 VDD.t2127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X199 VDD.t2126 a_7847_3425.t4 a_7752_3410.t1 VDD.t2125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X200 a_742_3184.t1 RWLB[2].t0 a_290_n953.t45 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X201 VSS.t2279 a_947_2421.t3 a_852_2406.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X202 a_7765_n953.t37 RWL[6].t0 a_7765_2180.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 a_1743_n2086.t0 a_1502_n2234.t2 VSS.t802 VSS.t801 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X204 a_6615_n953.t16 VSS.t751 a_6615_4148.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 VSS.t901 a_1522_2943.t3 a_1892_2943.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 a_9613_n4470.t1 Iref0.t0 a_9672_n4114.t1 VSS.t2232 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X207 VDD.t2098 a_372_3425.t3 a_277_3410.t1 VDD.t2097 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X208 a_2590_3666.t0 a_2577_3651.t3 VSS.t860 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X209 a_7283_n953.t8 WWLD[4].t2 a_7272_n271.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X210 VDD.t2096 a_n1233_n4483.t3 ADC2_OUT[0].t1 VDD.t2095 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X211 a_8020_4887.t20 PRE_SRAM.t0 VDD.t2012 VDD.t2011 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X212 a_4972_3666.t1 a_4877_3651.t3 VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_2097_1216.t2 a_2002_1201.t3 VDD.t468 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X214 VDD.t548 a_7847_452.t3 a_7752_437.t1 VDD.t547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X215 a_8217_n812.t0 VSS.t750 a_7765_n953.t2 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X216 a_1892_975.t1 RWLB[11].t1 a_1440_n953.t44 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X217 a_8433_n953.t2 WWL[11].t1 a_8422_975.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 VSS.t474 a_5547_3184.t3 a_5917_3184.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X219 a_545_4887.t22 PRE_SRAM.t1 VDD.t2014 VDD.t2013 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 VDD.t2207 a_4397_4445.t4 a_4302_4430.t1 VDD.t2206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X221 a_7283_n953.t0 WWL[1].t4 a_7272_3425.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 a_6615_3907.t1 a_6602_3892.t3 VSS.t856 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X223 a_958_n953.t26 WWL[11].t2 a_947_975.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 VDD.t95 PRE_CLSA.t4 ADC11_OUT[2].t0 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X225 VSS.t858 a_3247_4148.t3 a_3152_4133.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X226 VSS.t855 a_4397_2180.t3 a_4302_2165.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X227 VDD.t97 PRE_CLSA.t5 ADC8_OUT[2].t0 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X228 VDD.t2016 PRE_SRAM.t2 a_2108_n953.t3 VDD.t2015 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 VSS.t1042 a_8422_4445.t3 a_8792_4445.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X230 a_5917_693.t1 RWLB[12].t0 a_5465_n953.t20 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 a_8915_2943.t1 a_8902_2928.t3 VSS.t1548 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X232 a_3740_1939.t0 a_3727_1924.t3 VSS.t1550 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X233 a_6122_1939.t2 a_6027_1924.t3 VDD.t1283 VDD.t1282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X234 VSS.t1498 a_5632_n6430# a_6812_n6503.t1 VSS.t378 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X235 a_7847_3907.t2 a_7752_3892.t3 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X236 a_3165_3425.t1 a_3152_3410.t3 VSS.t1534 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 a_4618_n2086.t0 a_4377_n2234.t2 VSS.t973 VSS.t972 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 a_12963_n8583.t1 ADC14_OUT[3].t3 VDD.t1295 VDD.t1294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X239 a_4570_4887.t20 PRE_SRAM.t3 a_4408_n953.t22 VDD.t2017 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X240 a_372_2421.t1 a_277_2406.t3 VSS.t1062 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X241 VSS.t1061 a_947_1939.t3 a_1317_1939.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X242 a_7642_211.t0 RWLB[14].t0 a_7190_n953.t37 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 a_6122_693.t1 a_6027_678.t3 VSS.t1041 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X244 a_372_n271.t2 a_277_n286.t3 VSS.t2521 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X245 a_13171_n4470.t0 VCLP.t5 a_13033_n4470.t1 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X246 VDD.t1285 a_1522_452.t3 a_1427_437.t0 VDD.t1284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X247 a_7302_n1770.t1 a_7283_n953.t27 a_7260_n1770.t2 VSS.t2295 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X248 a_7067_n512.t0 VSS.t749 a_6615_n953.t12 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X249 a_852_n527.t0 WWLD[5].t0 a_1120_4887.t4 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X250 VDD.t99 PRE_CLSA.t6 ADC1_OUT[2].t0 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X251 VDD.t1155 PRE_VLSA.t6 a_8935_n1371.t0 VDD.t1154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X252 a_7858_n953.t22 WWLD[0].t1 a_7847_4686.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 a_4397_3907.t0 a_4302_3892.t3 VSS.t1214 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X254 a_1522_1457.t0 a_1427_1442.t3 VSS.t1201 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X255 a_7190_n953.t14 VSS.t748 a_7190_4148.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X256 a_8422_3666.t1 a_8327_3651.t3 VDD.t910 VDD.t909 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X257 a_n2415_n5850.t0 PRE_CLSA.t7 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X258 VDD.t1990 a_2097_3184.t4 a_2002_3169.t1 VDD.t1989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X259 a_6697_2943.t1 a_6602_2928.t3 VSS.t462 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X260 a_1317_1698.t1 RWLB[8].t0 a_865_n953.t30 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 VSS.t1013 a_6122_693.t3 a_6492_693.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X262 a_3493_n5850.t1 ADC6_OUT[1].t3 a_3563_n5338.t2 VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X263 VSS.t1199 a_4972_n30.t3 a_4877_n45.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X264 a_2015_n953.t48 RWL[14].t1 a_2015_211.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X265 VDD.t1194 PRE_A.t0 a_5543_n2422.t1 VDD.t1193 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X266 a_1522_975.t2 a_1427_960.t3 VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X267 a_9178_n6503.t2 a_5743_n6391# a_9143_n6849.t1 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X268 VSS.t1491 a_6122_3184.t3 a_6492_3184.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X269 a_4302_2406.t1 WWL[5].t0 a_4570_4887.t4 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X270 a_7272_452.t2 a_7177_437.t3 VDD.t728 VDD.t727 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X271 VSS.t2240 a_947_211.t3 a_852_196.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X272 VDD.t2019 PRE_SRAM.t4 a_5558_n953.t4 VDD.t2018 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X273 a_7190_3907.t1 a_7177_3892.t3 VSS.t2195 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X274 a_6615_3425.t1 a_6602_3410.t3 VSS.t89 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X275 a_8340_n953.t47 RWL[5].t1 a_8340_2421.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X276 a_7765_1457.t1 a_7752_1442.t3 VSS.t1300 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X277 a_4302_n286.t1 WWLD[4].t3 a_4570_4887.t16 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X278 a_4883_n8071.t1 Iref3.t1 a_4942_n8026.t1 VSS.t1981 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X279 VSS.t1090 a_3822_4148.t3 a_3727_4133.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X280 a_3740_n953.t47 RWL[14].t2 a_3740_211.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X281 a_n279_n6503.t2 a_n52_n7216.t3 ADC3_OUT[2].t1 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X282 a_865_n953.t45 RWL[5].t2 a_865_2421.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X283 VDD.t1394 a_8997_4686.t4 a_8902_4671.t1 VDD.t1393 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X284 a_7847_3425.t2 a_7752_3410.t3 VDD.t1966 VDD.t1965 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 VSS.t1069 a_4397_2421.t3 a_4767_2421.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X286 VSS.t1546 a_2672_211.t3 a_2577_196.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X287 a_383_n953.t11 WWLD[5].t1 a_372_n512.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X288 a_7247_n8071.t1 Iref3.t2 a_7306_n8026.t1 VSS.t1982 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X289 a_8221_n8583.t2 PRE_CLSA.t8 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X290 VDD.t1196 PRE_A.t1 a_3231_n4378.t3 VDD.t1195 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X291 a_6602_4133.t0 WWLD[2].t0 a_6870_4887.t15 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X292 VSS.t466 a_6697_2943.t3 a_7067_2943.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X293 a_7847_3907.t1 a_7752_3892.t4 VSS.t81 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X294 a_2097_4445.t1 a_2002_4430.t3 VDD.t708 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X295 a_1440_n953.t7 VSS.t747 a_1440_3907.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X296 VSS.t1517 a_4972_2421.t3 a_4877_2406.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X297 VDD.t692 a_2672_4148.t3 a_2577_4133.t2 VDD.t691 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 VDD.t410 a_5547_3184.t4 a_5452_3169.t0 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X299 VDD.t361 a_3822_2180.t3 a_3727_2165.t1 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X300 a_4972_1939.t1 a_4877_1924.t3 VSS.t50 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X301 VSS.t2030 a_372_452.t3 a_742_452.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X302 VSS.t267 SAEN.t2 a_13637_n3770.t0 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X303 a_4397_3425.t1 a_4302_3410.t3 VSS.t1790 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X304 a_8452_n1770.t1 a_8433_n953.t27 a_8410_n1770.t1 VSS.t2271 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X305 a_2590_n953.t17 VSS.t746 a_2590_n1053.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X306 VDD.t1802 a_3247_452.t3 a_3152_437.t1 VDD.t1801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 VDD.t105 PRE_CLSA.t9 ADC0_OUT[2].t0 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X308 a_1317_1216.t0 RWLB[10].t0 a_865_n953.t36 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X309 a_6027_n827.t0 WWLD[6].t0 a_6295_4887.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X310 a_8902_196.t1 WWL[14].t1 a_9170_4887.t19 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X311 a_n3792_n8026.t0 VCLP.t6 a_n3827_n7825.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X312 a_n3565_n5850.t0 PRE_CLSA.t10 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X313 a_11776_n4483.t0 PRE_CLSA.t11 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X314 a_11549_n3770.t1 a_11776_n4483.t3 ADC13_OUT[0].t2 VSS.t1856 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X315 VSS.t1101 a_8422_2180.t3 a_8327_2165.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X316 a_3165_n953.t35 RWL[8].t0 a_3165_1698.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 a_6122_1698.t1 a_6027_1683.t3 VSS.t2124 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X318 a_290_n30.t1 a_277_n45.t3 VSS.t435 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X319 VDD.t1198 PRE_A.t2 a_6693_n2422.t3 VDD.t1197 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X320 VSS.t1102 a_7272_4148.t3 a_7177_4133.t0 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X321 a_2015_n953.t24 RWL[0].t1 a_2015_3666.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X322 a_1317_211.t0 RWLB[14].t1 a_865_n953.t37 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 a_n3357_n4470.t0 VCLP.t7 a_n3495_n4470.t1 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X324 VDD.t2021 PRE_SRAM.t5 a_6133_n953.t21 VDD.t2020 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X325 a_4983_n953.t3 WWL[2].t2 a_4972_3184.t1 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X326 a_2519_n5338.t0 VCLP.t8 a_2381_n5338.t1 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X327 a_7190_3425.t0 a_7177_3410.t3 VSS.t1641 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X328 VDD.t1413 a_947_1939.t4 a_852_1924.t1 VDD.t1412 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 a_8997_452.t2 a_8902_437.t3 VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X330 a_3165_n953.t0 VSS.t745 a_3165_n812.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X331 VSS.t781 a_5118_n2426.t4 a_5595_n5092.t1 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X332 a_n1233_n4483.t1 ADC2_OUT[0].t3 a_n1163_n4470.t2 VSS.t900 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X333 a_8595_4887.t21 PRE_SRAM.t6 a_8433_n953.t4 VDD.t2022 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X334 a_8902_2647.t0 WWL[4].t0 a_9170_4887.t12 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 VSS.t1792 a_4972_1939.t3 a_5342_1939.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X336 a_1440_n953.t11 VSS.t744 a_1440_n271.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X337 a_n2345_n5338.t0 SAEN.t3 a_n2148_n5293.t0 VSS.t268 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X338 a_1522_4686.t1 a_1427_4671.t3 VSS.t777 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X339 a_1522_693.t1 a_1427_678.t3 VSS.t1634 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X340 a_4315_n30.t1 a_4302_n45.t3 VSS.t423 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X341 VSS.t1637 a_8997_1939.t3 a_8902_1924.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X342 a_4675_n7216.t1 ADC7_OUT[2].t3 VDD.t1228 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X343 a_2660_n1770.t2 a_2845_4887.t27 a_2853_n1770.t1 VSS.t384 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X344 VDD.t452 a_4972_2662.t3 a_4877_2647.t1 VDD.t451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X345 a_n52_n7216.t1 ADC3_OUT[2].t3 VDD.t682 VDD.t681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X346 a_5558_n953.t18 WWL[3].t0 a_5547_2943.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X347 a_2590_n953.t19 RWL[9].t0 a_2590_1457.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X348 a_8997_1457.t0 a_8902_1442.t3 VSS.t2163 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X349 a_4877_960.t0 WWL[11].t3 a_5145_4887.t26 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X350 a_4877_n527.t2 WWLD[5].t2 a_5145_4887.t2 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X351 a_1440_n953.t22 RWL[1].t0 a_1440_3425.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X352 a_7847_3425.t1 a_7752_3410.t4 VSS.t2235 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X353 VSS.t2516 a_927_n2234.t2 a_1050_n2132.t0 VSS.t2515 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X354 VSS.t1977 a_8997_2662.t3 a_9367_2662.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X355 a_5342_1698.t1 RWLB[8].t1 a_4890_n953.t39 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X356 VSS.t1294 a_1522_693.t3 a_1892_693.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X357 a_n2642_n5293.t2 a_n2415_n5850.t3 ADC1_OUT[1].t1 VSS.t1676 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X358 a_3042_452.t0 RWLB[13].t0 a_2590_n953.t22 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X359 a_7765_4686.t1 a_7752_4671.t3 VSS.t834 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 a_4408_n953.t19 WWL[6].t0 a_4397_2180.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X361 a_6615_n953.t37 RWL[8].t1 a_6615_1698.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X362 a_10797_n4470.t1 Iref0.t1 a_10856_n4114.t1 VSS.t2233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X363 a_2672_452.t1 a_2577_437.t3 VDD.t1738 VDD.t1737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X364 a_n2207_n7203.t1 Iref2.t0 a_n2148_n6847.t1 VSS.t1978 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X365 a_5630_n6503.t2 a_5857_n7216.t3 ADC8_OUT[2].t1 VSS.t1361 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X366 VSS.t270 SAEN.t4 a_6812_n3770.t0 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X367 a_3165_n953.t32 RWL[10].t2 a_3165_1216.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X368 a_6122_1216.t1 a_6027_1201.t3 VSS.t1609 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X369 VDD.t908 a_4397_2421.t4 a_4302_2406.t2 VDD.t907 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X370 a_5535_n1770.t2 a_5720_4887.t27 a_5728_n1770.t1 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X371 VSS.t2174 a_2672_n1053.t3 a_2577_n1068.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X372 a_6615_n953.t10 VSS.t743 a_6615_n812.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X373 a_5857_n4483.t2 ADC8_OUT[0].t3 VDD.t1550 VDD.t1549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X374 VDD.t394 a_n3565_n7216.t3 ADC0_OUT[2].t1 VDD.t362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X375 a_7994_n6503.t2 a_8221_n7216.t3 ADC10_OUT[2].t1 VSS.t243 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X376 a_1522_2180.t2 a_1427_2165.t3 VDD.t1386 VDD.t1385 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X377 VDD.t111 PRE_CLSA.t12 ADC12_OUT[2].t0 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X378 VSS.t845 a_3802_n2234.t2 a_3925_n2132.t0 VSS.t844 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 VSS.t822 a_8422_2421.t3 a_8792_2421.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X380 VSS.t1649 a_3247_1698.t3 a_3152_1683.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X381 VDD.t113 PRE_CLSA.t13 ADC4_OUT[0].t0 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X382 a_3833_n953.t17 WWL[7].t2 a_3822_1939.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X383 a_8217_975.t0 RWLB[11].t2 a_7765_n953.t24 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X384 a_8327_n527.t2 WWLD[5].t3 a_8595_4887.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X385 a_1317_4445.t0 VSS.t742 a_865_n953.t18 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X386 VDD.t1904 a_6697_4148.t3 a_6602_4133.t1 VDD.t1903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 VSS.t960 a_3247_n812.t3 a_3152_n827.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X388 a_9178_n3770.t1 VCLP.t9 a_9143_n4116.t0 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X389 VSS.t1788 a_1522_3907.t3 a_1892_3907.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X390 a_5342_1216.t0 RWLB[10].t1 a_4890_n953.t45 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X391 VSS.t957 a_2077_n2234.t2 a_2200_n2132.t0 VSS.t956 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X392 a_2002_3651.t2 WWL[0].t2 a_2270_4887.t22 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 a_7858_n953.t16 WWL[4].t1 a_7847_2662.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X394 a_4302_196.t1 WWL[14].t2 a_4570_4887.t17 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 VDD.t1758 a_7847_n30.t3 a_7752_n45.t2 VDD.t1757 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X396 a_5465_n953.t12 VSS.t741 a_5465_n512.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X397 a_6040_n953.t27 RWL[0].t2 a_6040_3666.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X398 a_7190_n953.t29 RWL[8].t2 a_7190_1698.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X399 VSS.t1298 a_2672_1457.t3 a_2577_1442.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X400 a_6615_n953.t35 RWL[10].t3 a_6615_1216.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X401 a_n279_n3770.t2 a_n52_n4483.t3 ADC3_OUT[0].t2 VSS.t1251 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X402 VDD.t1730 a_8422_1939.t3 a_8327_1924.t2 VDD.t1729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X403 a_13171_n4470.t1 Iref0.t2 a_13230_n4114.t1 VSS.t2234 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X404 a_9367_1939.t1 RWLB[7].t0 a_8915_n953.t38 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X405 a_4397_452.t2 a_4302_437.t3 VDD.t952 VDD.t951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X406 a_7190_n953.t18 VSS.t740 a_7190_n812.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X407 VSS.t1989 a_2097_3666.t3 a_2467_3666.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X408 a_4192_n30.t0 RWLB[15].t0 a_3740_n953.t35 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X409 a_4890_3184.t1 a_4877_3169.t3 VSS.t438 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X410 a_3152_1924.t2 WWL[7].t3 a_3420_4887.t17 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X411 a_958_n953.t15 WWL[15].t0 a_947_n30.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X412 VSS.t1605 a_2097_n512.t3 a_2002_n527.t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X413 a_2590_n953.t11 VSS.t739 a_2590_4686.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X414 a_8997_4686.t1 a_8902_4671.t3 VSS.t2502 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X415 a_947_4148.t1 a_852_4133.t3 VDD.t1752 VDD.t1751 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X416 a_7272_3184.t2 a_7177_3169.t3 VDD.t1185 VDD.t1184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X417 VDD.t1153 PRE_VLSA.t7 a_310_n1371.t0 VDD.t1152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X418 VSS.t1311 a_3822_1698.t3 a_3727_1683.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X419 VDD.t1552 a_8997_2662.t4 a_8902_2647.t1 VDD.t1551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 VSS.t1986 a_3247_1216.t3 a_3152_1201.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X421 a_277_678.t2 WWL[12].t3 a_545_4887.t7 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X422 VSS.t436 a_8997_452.t3 a_8902_437.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X423 VDD.t1998 a_3493_n8583.t3 ADC6_OUT[3].t2 VDD.t1997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X424 VSS.t1246 a_4952_n2234.t2 a_5075_n2132.t0 VSS.t1245 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X425 a_2097_975.t0 a_2002_960.t3 VSS.t879 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X426 VSS.t1778 a_1522_n271.t3 a_1892_n271.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X427 VSS.t2182 a_3822_n812.t3 a_3727_n827.t2 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X428 a_1440_n812.t1 a_1427_n827.t3 VSS.t877 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X429 a_2097_2421.t1 a_2002_2406.t3 VDD.t1705 VDD.t1704 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X430 a_6602_1683.t2 WWL[8].t0 a_6870_4887.t5 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 a_6615_n953.t23 RWL[15].t0 a_6615_n30.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X432 a_8915_n953.t16 VSS.t738 a_8915_n512.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 a_5452_3651.t2 WWL[0].t3 a_5720_4887.t24 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X434 a_8433_n953.t25 WWL[6].t1 a_8422_2180.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 a_2178_n2086.t0 WE.t4 a_2108_n953.t12 VSS.t2407 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X436 a_3165_n953.t15 VSS.t737 a_3165_4445.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X437 a_6122_4445.t0 a_6027_4430.t3 VSS.t1323 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X438 a_742_3666.t0 RWLB[0].t0 a_290_n953.t25 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X439 a_2097_n271.t1 a_2002_n286.t3 VDD.t1898 VDD.t1897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X440 a_n52_n5850.t0 PRE_CLSA.t14 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X441 a_372_n1053.t1 a_277_n1068.t3 VDD.t822 VDD.t821 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X442 VSS.t1913 a_1522_3425.t3 a_1892_3425.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X443 VSS.t2104 a_6697_975.t3 a_6602_960.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X444 a_5558_n953.t9 WWL[12].t4 a_5547_693.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 a_13864_n5850.t1 ADC15_OUT[1].t4 a_13934_n5338.t2 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X446 a_958_n953.t16 WWL[6].t2 a_947_2180.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X447 VDD.t642 a_2672_1698.t3 a_2577_1683.t1 VDD.t641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X448 VSS.t2450 a_7847_n1053.t3 a_7752_n1068.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X449 a_4315_2180.t0 a_4302_2165.t3 VSS.t477 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X450 a_7190_n953.t2 RWL[10].t4 a_7190_1216.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X451 a_6027_196.t2 WWL[14].t3 a_6295_4887.t16 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X452 a_7283_n953.t10 WWL[14].t4 a_7272_211.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X453 VSS.t1656 a_5547_3666.t3 a_5917_3666.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_7847_693.t0 a_7752_678.t3 VSS.t1346 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X455 a_4883_n5338.t0 VCLP.t10 a_4745_n5338.t1 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X456 VDD.t1396 a_2672_n812.t3 a_2577_n827.t2 VDD.t1395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X457 a_4397_4148.t2 a_4302_4133.t3 VDD.t1573 VDD.t1572 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X458 a_5547_2180.t2 a_5452_2165.t3 VDD.t1859 VDD.t1858 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 a_3727_1442.t2 WWL[9].t2 a_3995_4887.t23 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X460 VSS.t1148 a_5547_n512.t3 a_5452_n527.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X461 a_9008_n953.t7 WWL[7].t4 a_8997_1939.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X462 a_865_452.t0 a_852_437.t4 VSS.t2431 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X463 VSS.t424 a_7272_1698.t3 a_7177_1683.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X464 VSS.t1155 a_6268_n2426.t4 a_7959_n5092.t1 VSS.t1153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X465 a_8902_2928.t2 WWL[3].t1 a_9170_4887.t10 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X466 a_7247_n5338.t0 VCLP.t11 a_7109_n5338.t1 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X467 VSS.t1820 a_3822_1216.t3 a_3727_1201.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X468 a_3617_975.t0 RWLB[11].t3 a_3165_n953.t22 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X469 VSS.t2131 a_7418_n2426.t4 a_10327_n5092.t1 VSS.t2129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X470 a_9367_452.t0 RWLB[13].t1 a_8915_n953.t24 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X471 VSS.t1723 a_7272_n812.t3 a_7177_n827.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X472 a_5342_4445.t0 VSS.t736 a_4890_n953.t13 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X473 VSS.t2200 a_6697_3907.t3 a_7067_3907.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X474 a_1522_2662.t0 a_1427_2647.t3 VSS.t1665 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X475 a_2097_2180.t1 a_2002_2165.t4 VSS.t1273 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X476 a_8340_693.t0 a_8327_678.t3 VSS.t893 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X477 a_5547_n30.t2 a_5452_n45.t3 VDD.t1736 VDD.t1735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X478 a_5857_n4483.t0 PRE_CLSA.t15 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X479 VSS.t1776 a_2672_4686.t3 a_2577_4671.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X480 a_6615_n953.t5 VSS.t735 a_6615_4445.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 a_5630_n3770.t2 a_5857_n4483.t3 ADC8_OUT[0].t1 VSS.t1341 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X482 VSS.t2256 a_7847_1457.t3 a_7752_1442.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X483 a_6602_1201.t2 WWL[10].t1 a_6870_4887.t8 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X484 VDD.t1519 a_1522_n512.t3 a_1427_n527.t1 VDD.t1518 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 a_3328_n2086.t1 WE.t5 a_3258_n953.t5 VSS.t2408 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 a_947_n1053.t0 a_852_n1068.t3 VSS.t1965 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X487 a_383_n953.t24 WWLD[2].t1 a_372_4148.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 VDD.t1742 a_2097_3666.t4 a_2002_3651.t0 VDD.t1741 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X489 a_7765_2662.t1 a_7752_2647.t3 VSS.t1766 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 VDD.t528 a_2672_1216.t3 a_2577_1201.t2 VDD.t527 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X491 a_7994_n3770.t2 a_8221_n4483.t3 ADC10_OUT[0].t2 VSS.t874 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X492 a_10362_n6503.t0 a_10589_n7216.t3 ADC12_OUT[2].t1 VSS.t1564 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X493 VSS.t1727 a_3247_4445.t3 a_3152_4430.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X494 VDD.t1815 a_6677_n2234.t2 a_6800_n2132.t1 VDD.t1814 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X495 a_2672_n812.t1 a_2577_n827.t3 VSS.t1344 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X496 VSS.t2113 a_6122_3666.t3 a_6492_3666.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X497 a_7177_1924.t0 WWL[7].t5 a_7445_4887.t7 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X498 VSS.t1888 a_6122_n512.t3 a_6027_n527.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X499 a_3740_n512.t1 a_3727_n527.t3 VSS.t2374 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 a_5465_n953.t42 RWL[13].t0 a_5465_452.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X501 a_6122_n512.t2 a_6027_n527.t3 VDD.t1670 VDD.t1669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X502 a_3042_3184.t0 RWLB[2].t1 a_2590_n953.t48 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X503 VSS.t1456 a_7272_1216.t3 a_7177_1201.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X504 VSS.t1658 a_7847_693.t3 a_8217_693.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X505 a_10589_n4483.t2 ADC12_OUT[0].t3 VDD.t1452 VDD.t1451 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X506 VSS.t77 a_6697_n271.t4 a_7067_n271.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X507 a_n2415_n8583.t1 ADC1_OUT[3].t3 VDD.t1450 VDD.t1449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X508 VSS.t1166 a_4397_452.t3 a_4302_437.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X509 VDD.t1459 a_7272_n1053.t3 a_7177_n1068.t2 VDD.t1458 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X510 a_4315_n953.t46 RWL[2].t2 a_4315_3184.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X511 a_5547_2180.t1 a_5452_2165.t4 VSS.t1347 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X512 VSS.t2514 a_7847_975.t3 a_8217_975.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X513 VSS.t1702 a_372_211.t3 a_277_196.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X514 SA_OUT[0].t2 a_310_n1371.t3 a_553_n1770.t0 VSS.t1464 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X515 VSS.t2418 a_6697_3425.t4 a_7067_3425.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X516 VDD.t1677 a_7039_n5850.t3 ADC9_OUT[1].t1 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X517 a_5558_n953.t8 WWLD[3].t4 a_5547_3907.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X518 a_3258_n953.t26 WWL[11].t4 a_3247_975.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X519 a_593_n2086.t0 a_352_n2234.t2 VSS.t908 VSS.t907 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 a_372_n812.t2 a_277_n827.t3 VDD.t696 VDD.t695 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X521 a_7190_n953.t17 VSS.t734 a_7190_4445.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X522 a_1317_2421.t0 RWLB[5].t1 a_865_n953.t47 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X523 VDD.t694 a_6697_1698.t3 a_6602_1683.t0 VDD.t693 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 a_1317_n271.t0 VSS.t733 a_865_n953.t13 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X525 VSS.t1193 a_372_n1053.t3 a_742_n1053.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X526 a_1892_n812.t0 VSS.t732 a_1440_n953.t12 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 VDD.t1398 a_5547_3666.t4 a_5452_3651.t0 VDD.t1397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X528 a_3727_4671.t0 WWLD[0].t2 a_3995_4887.t7 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X529 a_8340_2180.t0 a_8327_2165.t3 VSS.t2122 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X530 VSS.t2077 a_947_3184.t3 a_852_3169.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X531 a_3247_211.t0 a_3152_196.t3 VSS.t1034 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X532 a_1427_196.t2 WWL[14].t5 a_1695_4887.t19 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X533 a_2683_n953.t9 WWL[14].t6 a_2672_211.t1 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X534 a_2108_n953.t7 WWLD[5].t4 a_2097_n512.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X535 a_2672_3907.t2 a_2577_3892.t3 VDD.t1664 VDD.t1663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 a_865_2180.t1 a_852_2165.t3 VSS.t1036 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X537 VDD.t1358 a_6697_n812.t3 a_6602_n827.t2 VDD.t1357 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 a_3740_n953.t41 RWL[3].t1 a_3740_2943.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 a_3493_n5850.t0 PRE_CLSA.t16 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X540 VSS.t1052 a_3822_4445.t3 a_3727_4430.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X541 a_4767_2180.t1 RWLB[6].t3 a_4315_n953.t38 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 a_2015_693.t0 a_2002_678.t3 VSS.t1884 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X543 a_3617_4148.t0 VSS.t731 a_3165_n953.t10 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X544 a_277_1442.t0 WWL[9].t3 a_545_4887.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X545 a_6602_960.t2 WWL[11].t5 a_6870_4887.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X546 a_902_n5293.t1 VCLP.t12 a_867_n5092.t0 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X547 a_3802_n2234.t0 Din[6].t0 VSS.t1615 VSS.t1614 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X548 a_4983_n953.t26 WWL[0].t4 a_4972_3666.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X549 VDD.t440 a_7272_1457.t3 a_7177_1442.t1 VDD.t439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X550 a_4972_211.t1 a_4877_196.t3 VSS.t505 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X551 VSS.t1672 a_7847_4686.t3 a_7752_4671.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X552 a_8997_2662.t0 a_8902_2647.t4 VSS.t2338 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X553 a_4767_452.t0 RWLB[13].t2 a_4315_n953.t22 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X554 a_6602_4430.t2 WWLD[1].t1 a_6870_4887.t25 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X555 a_2590_n953.t44 RWL[4].t1 a_2590_2662.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X556 a_742_211.t1 RWLB[14].t2 a_290_n953.t39 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X557 a_5558_n953.t13 WWLD[4].t4 a_5547_n271.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X558 a_8429_n5338.t1 Iref1.t1 a_8488_n5293.t1 VSS.t2220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X559 a_947_1698.t1 a_852_1683.t3 VDD.t1340 VDD.t1339 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X560 a_3740_693.t0 a_3727_678.t4 VSS.t248 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X561 a_6708_n953.t26 WWL[11].t6 a_6697_975.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X562 VSS.t1026 a_372_1457.t3 a_742_1457.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X563 a_2084_n8026.t2 a_2311_n8583.t3 ADC5_OUT[3].t0 VSS.t1106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X564 VDD.t594 a_2672_4445.t3 a_2577_4430.t1 VDD.t593 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X565 a_372_3184.t1 a_277_3169.t3 VSS.t1695 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X566 a_1129_n8583.t1 ADC4_OUT[3].t3 VDD.t666 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X567 a_4972_n512.t1 a_4877_n527.t3 VSS.t924 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X568 a_5558_n953.t0 WWL[1].t5 a_5547_3425.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X569 VSS.t1022 a_n2677_n4378.t4 a_n2677_n6849.t1 VSS.t1021 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X570 a_6677_n2234.t0 Din[11].t0 VSS.t993 VSS.t992 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X571 a_3165_n953.t46 RWL[5].t3 a_3165_2421.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X572 a_6122_2421.t0 a_6027_2406.t3 VSS.t1049 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X573 VDD.t652 a_6697_1216.t3 a_6602_1201.t1 VDD.t651 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X574 a_7039_n7216.t0 PRE_CLSA.t17 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X575 VDD.t592 a_2097_693.t3 a_2002_678.t0 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X576 a_6122_n271.t0 a_6027_n286.t3 VSS.t1031 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X577 VSS.t441 a_7272_4445.t3 a_7177_4430.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X578 a_372_452.t0 a_277_437.t3 VDD.t387 VDD.t386 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X579 a_8020_4887.t25 WE.t6 a_8068_n2086.t0 VSS.t2379 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X580 a_290_4148.t1 a_277_4133.t3 VSS.t1318 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X581 a_2672_3425.t2 a_2577_3410.t3 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X582 a_4192_4148.t1 VSS.t730 a_3740_n953.t18 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X583 VDD.t2283 a_7847_975.t4 a_7752_960.t1 VDD.t2282 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X584 a_2381_n8071.t1 SAEN.t5 a_2578_n8026.t0 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X585 VSS.t1831 a_3247_693.t3 a_3617_693.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 a_n2207_n8071.t0 VCLP.t13 a_n2345_n8071.t1 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X587 VDD.t123 PRE_CLSA.t18 ADC7_OUT[3].t0 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X588 a_4302_3169.t0 WWL[2].t3 a_4570_4887.t22 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X589 a_3277_n1770.t0 a_3258_n953.t27 a_3235_n1770.t1 VSS.t2419 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X590 a_4397_1698.t2 a_4302_1683.t3 VDD.t2150 VDD.t2149 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X591 VDD.t1334 a_372_975.t3 a_277_960.t2 VDD.t1333 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X592 a_4952_n2234.t0 Din[8].t0 VSS.t1223 VSS.t1222 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X593 a_5465_n953.t11 VSS.t729 a_5465_4148.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X594 a_8422_4148.t1 a_8327_4133.t3 VSS.t1226 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X595 a_8340_n953.t0 RWL[2].t3 a_8340_3184.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X596 a_8327_960.t2 WWL[11].t7 a_8595_4887.t26 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 a_n1233_n4483.t0 PRE_CLSA.t19 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X598 VSS.t1619 a_4972_211.t3 a_5342_211.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X599 VDD.t1336 a_13864_n8583.t3 ADC15_OUT[3].t1 VDD.t1335 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X600 a_947_4148.t0 a_852_4133.t4 VSS.t1992 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X601 a_865_n953.t0 RWL[2].t4 a_865_3184.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X602 a_1522_2943.t2 a_1427_2928.t3 VSS.t1886 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X603 a_947_1216.t2 a_852_1201.t3 VDD.t1232 VDD.t1231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X604 VDD.t1654 a_1129_n4483.t3 ADC4_OUT[0].t1 VDD.t1653 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X605 a_2015_n1053.t1 a_2002_n1068.t3 VSS.t895 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 a_7067_n812.t1 VSS.t728 a_6615_n953.t14 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X607 a_5342_2421.t0 RWLB[5].t2 a_4890_n953.t22 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X608 a_7283_n953.t1 WWL[11].t8 a_7272_975.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X609 a_852_n827.t0 WWLD[6].t1 a_1120_4887.t13 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X610 VSS.t1905 a_4397_3184.t3 a_4767_3184.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X611 a_5342_n271.t0 VSS.t727 a_4890_n953.t14 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X612 a_5465_3907.t1 a_5452_3892.t3 VSS.t1830 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X613 VSS.t813 a_2672_2662.t3 a_2577_2647.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X614 a_6615_n953.t47 RWL[5].t4 a_6615_2421.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X615 VDD.t127 PRE_CLSA.t20 ADC2_OUT[3].t0 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X616 VSS.t386 a_2097_4148.t3 a_2002_4133.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X617 VSS.t1514 a_4972_3184.t3 a_4877_3169.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X618 a_10362_n3770.t2 a_10589_n4483.t3 ADC12_OUT[0].t1 VSS.t1815 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X619 a_8985_n1770.t0 PRE_VLSA.t8 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X620 a_1552_n1770.t0 a_1533_n953.t27 a_1510_n1770.t0 VSS.t897 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X621 a_2590_1939.t1 a_2577_1924.t3 VSS.t1834 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 a_6133_n953.t4 WWLD[5].t5 a_6122_n512.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X623 a_277_4671.t1 WWLD[0].t3 a_545_4887.t21 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_7765_2943.t1 a_7752_2928.t3 VSS.t1853 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X625 a_4972_1939.t2 a_4877_1924.t4 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X626 VDD.t570 a_7272_4686.t3 a_7177_4671.t2 VDD.t569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X627 a_7827_n2234.t0 Din[13].t0 VSS.t1486 VSS.t1485 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X628 a_7642_4148.t0 VSS.t726 a_7190_n953.t6 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X629 a_8792_2180.t1 RWLB[6].t4 a_8340_n953.t38 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X630 a_2577_2165.t0 WWL[6].t3 a_2845_4887.t12 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 a_383_n953.t23 WWL[8].t1 a_372_1698.t1 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X632 VSS.t272 SAEN.t6 a_n3792_n6503.t0 VSS.t262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X633 a_9170_4887.t7 WE.t7 a_9218_n2086.t1 VSS.t2380 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X634 a_1427_4133.t0 WWLD[2].t2 a_1695_4887.t17 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X635 a_8915_n953.t14 VSS.t725 a_8915_4148.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X636 VSS.t1839 a_3247_2421.t3 a_3152_2406.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X637 a_12963_n5850.t1 ADC14_OUT[1].t3 VDD.t1238 VDD.t1237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X638 VSS.t1007 a_372_4686.t3 a_742_4686.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X639 a_n279_n6503.t1 VCLP.t14 a_n314_n6849.t0 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X640 a_4890_3666.t0 a_4877_3651.t4 VSS.t472 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X641 a_383_n953.t17 WWLD[6].t2 a_372_n812.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X642 a_7272_3666.t1 a_7177_3651.t3 VDD.t2152 VDD.t2151 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X643 a_7283_n953.t19 WWL[15].t1 a_7272_n30.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X644 a_8221_n7216.t2 ADC10_OUT[2].t4 a_8291_n7203.t0 VSS.t246 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X645 a_4397_1216.t1 a_4302_1201.t3 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X646 a_4427_n1770.t1 a_4408_n953.t27 a_4385_n1770.t1 VSS.t2304 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X647 a_8402_n2234.t1 Din[14].t0 VDD.t636 VDD.t635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X648 VDD.t1465 a_6697_4445.t3 a_6602_4430.t0 VDD.t1464 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X649 VSS.t1709 a_6122_n30.t3 a_6492_n30.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X650 a_8915_3907.t1 a_8902_3892.t3 VSS.t1290 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X651 VSS.t47 a_6697_2180.t3 a_6602_2165.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X652 VSS.t935 a_5547_4148.t3 a_5452_4133.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X653 VDD.t2024 PRE_SRAM.t7 a_4408_n953.t23 VDD.t2023 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X654 a_5465_3425.t1 a_5452_3410.t3 VSS.t1746 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X655 a_7190_n953.t47 RWL[5].t5 a_7190_2421.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X656 a_8422_1939.t2 a_8327_1924.t3 VDD.t1964 VDD.t1963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X657 a_6870_4887.t4 PRE_SRAM.t8 a_6708_n953.t22 VDD.t2025 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X658 VSS.t1316 a_3247_1939.t3 a_3617_1939.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 a_3727_2647.t2 WWL[4].t2 a_3995_4887.t24 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X660 a_7642_n30.t1 RWLB[15].t1 a_7190_n953.t33 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X661 a_7752_437.t2 WWL[13].t1 a_8020_4887.t19 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X662 a_9367_n512.t0 VSS.t724 a_8915_n953.t3 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X663 a_383_n953.t7 WWL[10].t2 a_372_1216.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X664 a_3266_n5293.t2 VCLP.t15 a_3231_n5092.t0 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X665 a_6697_3907.t0 a_6602_3892.t4 VSS.t857 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X666 VSS.t872 a_3822_2421.t3 a_3727_2406.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X667 a_3152_n527.t0 WWLD[5].t6 a_3420_4887.t13 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X668 a_947_4445.t2 a_852_4430.t3 VDD.t2193 VDD.t2192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 a_3822_1457.t0 a_3727_1442.t3 VSS.t2136 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X670 a_5547_975.t1 a_5452_960.t3 VSS.t1434 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X671 a_3247_693.t1 a_3152_678.t3 VDD.t458 VDD.t457 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X672 a_8221_n5850.t0 PRE_CLSA.t21 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X673 VDD.t1043 a_1522_4148.t3 a_1427_4133.t1 VDD.t1042 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X674 VDD.t1681 a_4397_3184.t4 a_4302_3169.t1 VDD.t1680 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X675 a_8997_2943.t1 a_8902_2928.t4 VSS.t1549 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X676 a_3617_1698.t1 RWLB[8].t2 a_3165_n953.t36 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X677 VSS.t1436 a_6697_n30.t3 a_6602_n45.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X678 VSS.t274 SAEN.t7 a_12736_n8026.t0 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X679 VSS.t234 a_8422_3184.t3 a_8792_3184.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X680 VSS.t1797 a_7847_2662.t3 a_7752_2647.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X681 a_9008_n953.t8 WWL[14].t7 a_8997_211.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X682 a_9405_n8583.t0 PRE_CLSA.t22 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X683 VSS.t95 a_n3827_n4378.t0 a_n3827_n4378.t1 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X684 a_4877_n827.t2 WWLD[6].t3 a_5145_4887.t6 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X685 VDD.t2027 PRE_SRAM.t9 a_7858_n953.t24 VDD.t2026 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X686 a_6602_2406.t2 WWL[5].t1 a_6870_4887.t11 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X687 VDD.t1041 a_8422_693.t3 a_8327_678.t2 VDD.t1040 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X688 a_4448_n8026.t2 a_4675_n8583.t3 ADC7_OUT[3].t1 VSS.t1449 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X689 VSS.t98 a_4393_n2422.t0 a_4393_n2422.t1 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X690 a_6602_n286.t2 WWLD[4].t5 a_6870_4887.t14 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X691 a_8915_3425.t1 a_8902_3410.t3 VSS.t1430 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X692 VSS.t2463 a_6122_4148.t3 a_6027_4133.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X693 VDD.t550 a_2672_2421.t3 a_2577_2406.t1 VDD.t549 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X694 a_8997_1457.t1 a_8902_1442.t4 VDD.t1910 VDD.t1909 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X695 a_6040_975.t0 a_6027_960.t4 VSS.t2526 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X696 VSS.t1437 a_6697_n30.t4 a_7067_n30.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X697 VDD.t560 a_4972_2943.t3 a_4877_2928.t2 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X698 a_290_n953.t23 RWL[7].t0 a_290_1939.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X699 a_2590_n953.t23 RWL[15].t1 a_2590_n30.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X700 a_7752_2165.t0 WWL[6].t4 a_8020_4887.t12 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X701 VSS.t1410 a_8997_2943.t3 a_9367_2943.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X702 VSS.t951 a_3822_1939.t3 a_4192_1939.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X703 a_3740_n953.t11 VSS.t723 a_3740_3907.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X704 VSS.t2375 a_7272_2421.t3 a_7177_2406.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X705 a_4745_n8071.t0 SAEN.t8 a_4942_n8026.t0 VSS.t275 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X706 a_4397_4445.t2 a_4302_4430.t3 VDD.t2197 VDD.t2196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X707 a_1440_n953.t23 RWL[11].t0 a_1440_975.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X708 a_6697_3425.t0 a_6602_3410.t4 VSS.t83 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X709 VSS.t1669 a_7847_2180.t3 a_8217_2180.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X710 a_290_1698.t1 a_277_1683.t3 VSS.t1668 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X711 a_n3565_n8583.t1 ADC0_OUT[3].t3 a_n3495_n8071.t2 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X712 a_4890_n953.t7 VSS.t722 a_4890_n1053.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X713 a_4192_1698.t1 RWLB[8].t3 a_3740_n953.t32 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X714 a_3042_3666.t0 RWLB[0].t1 a_2590_n953.t25 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X715 a_3617_1216.t0 RWLB[10].t2 a_3165_n953.t40 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X716 a_7109_n8071.t0 SAEN.t9 a_7306_n8026.t0 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X717 VDD.t1400 SA_OUT[8].t3 a_4910_n1371.t1 VDD.t1399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X718 a_8327_n827.t0 WWLD[6].t4 a_8595_4887.t8 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X719 a_8902_n45.t2 WWL[15].t2 a_9170_4887.t14 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X720 a_2108_n953.t24 WWLD[2].t3 a_2097_4148.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X721 a_3258_n953.t13 WWL[6].t5 a_3247_2180.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X722 a_4315_n953.t47 RWL[0].t3 a_4315_3666.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X723 a_5465_n953.t33 RWL[8].t3 a_5465_1698.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X724 a_8422_1698.t1 a_8327_1683.t3 VSS.t1038 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X725 a_6812_n8026.t1 VCLP.t16 a_6777_n7825.t0 VSS.t178 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X726 VDD.t2029 PRE_SRAM.t10 a_8433_n953.t3 VDD.t2028 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X727 a_1317_n30.t1 RWLB[15].t2 a_865_n953.t34 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X728 VDD.t956 a_3247_1939.t4 a_3152_1924.t0 VDD.t955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X729 a_947_1698.t0 a_852_1683.t4 VSS.t1590 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X730 VSS.t2427 a_1522_n1053.t3 a_1427_n1068.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X731 a_5465_n953.t9 VSS.t721 a_5465_n812.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X732 VSS.t278 SAEN.t10 a_n3792_n3770.t0 VSS.t277 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X733 a_383_n953.t25 WWLD[1].t2 a_372_4445.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X734 VSS.t2049 a_7272_1939.t3 a_7642_1939.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X735 a_3740_n953.t21 VSS.t720 a_3740_n271.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X736 a_3822_4686.t1 a_3727_4671.t3 VSS.t1601 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X737 a_2097_3184.t2 a_2002_3169.t3 VDD.t2002 VDD.t2001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X738 VSS.t1210 a_5543_n2422.t4 a_6777_n6849.t1 VSS.t1209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X739 a_7302_n1770.t0 SA_OUT[12].t3 a_7210_n1371.t1 VSS.t2177 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X740 VDD.t337 SA_OUT[5].t3 a_3185_n1371.t2 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X741 VSS.t2478 a_2097_1698.t3 a_2002_1683.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X742 a_3152_437.t2 WWL[13].t2 a_3420_4887.t19 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X743 a_5465_211.t1 a_5452_196.t4 VSS.t160 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X744 a_3165_n953.t21 RWL[15].t2 a_3165_n30.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X745 a_n279_n3770.t1 VCLP.t17 a_n314_n4116.t0 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X746 VSS.t1393 a_947_3666.t3 a_852_3651.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X747 a_277_2647.t2 WWL[4].t3 a_545_4887.t15 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X748 VDD.t351 a_7272_2662.t3 a_7177_2647.t1 VDD.t350 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X749 a_8915_n953.t48 RWL[13].t1 a_8915_452.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X750 a_383_n953.t15 WWL[14].t8 a_372_211.t1 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X751 a_7858_n953.t13 WWL[3].t2 a_7847_2943.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X752 a_2683_n953.t8 WWL[7].t6 a_2672_1939.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X753 a_947_693.t1 a_852_678.t3 VSS.t2269 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X754 a_8291_n5338.t0 SAEN.t11 a_8488_n5293.t0 VSS.t279 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X755 a_8221_n4483.t1 ADC10_OUT[0].t3 a_8291_n4470.t2 VSS.t1698 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X756 a_7177_n527.t0 WWLD[5].t7 a_7445_4887.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X757 a_3740_n953.t24 RWL[1].t1 a_3740_3425.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X758 a_4890_n953.t18 RWL[9].t1 a_4890_1457.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X759 VSS.t468 a_372_1939.t3 a_277_1924.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X760 VSS.t459 a_2097_n812.t3 a_2002_n827.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X761 a_7642_1698.t1 RWLB[8].t4 a_7190_n953.t30 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X762 a_6697_452.t2 a_6602_437.t3 VSS.t1802 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X763 VSS.t232 a_2672_n30.t4 a_2577_n45.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X764 a_290_1216.t1 a_277_1201.t4 VSS.t390 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X765 a_9178_n6503.t1 a_9405_n7216.t4 ADC11_OUT[2].t1 VSS.t1440 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X766 a_6708_n953.t18 WWL[6].t6 a_6697_2180.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X767 a_1427_1683.t0 WWL[8].t2 a_1695_4887.t21 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X768 a_2311_n4483.t0 PRE_CLSA.t23 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X769 VSS.t906 a_372_2662.t3 a_742_2662.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X770 a_8915_n953.t19 RWL[8].t4 a_8915_1698.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X771 a_8997_4686.t2 a_8902_4671.t4 VDD.t2285 VDD.t2284 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X772 a_4192_1216.t1 RWLB[10].t3 a_3740_n953.t37 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X773 a_4408_n953.t11 WWL[14].t9 a_4397_211.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X774 a_5577_n1770.t1 SA_OUT[9].t3 a_5485_n1371.t1 VSS.t1432 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X775 SA_OUT[0].t0 PRE_VLSA.t9 VDD.t1151 VDD.t1150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X776 a_7765_n1053.t1 a_7752_n1068.t3 VSS.t1160 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X777 VDD.t85 a_3822_693.t3 a_3727_678.t0 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X778 a_9405_n4483.t1 ADC11_OUT[0].t3 VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X779 VDD.t31 SA_OUT[10].t3 a_6060_n1371.t2 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X780 VSS.t1203 a_1522_1457.t3 a_1427_1442.t0 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X781 a_5465_n953.t31 RWL[10].t5 a_5465_1216.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X782 a_8422_1216.t0 a_8327_1201.t3 VSS.t503 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X783 VSS.t239 a_2672_n30.t5 a_3042_n30.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X784 a_8915_n953.t11 VSS.t719 a_8915_n812.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X785 VDD.t434 a_6697_2421.t3 a_6602_2406.t0 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X786 a_1440_975.t1 a_1427_960.t4 VSS.t967 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X787 a_8429_n7203.t1 Iref2.t1 a_8488_n6847.t1 VSS.t1979 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X788 a_372_3666.t1 a_277_3651.t3 VSS.t2202 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X789 VDD.t1039 a_8997_2943.t4 a_8902_2928.t0 VDD.t1038 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X790 a_8217_1457.t0 RWLB[9].t0 a_7765_n953.t39 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X791 a_947_1216.t1 a_852_1201.t4 VSS.t1477 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X792 a_7190_452.t1 a_7177_437.t4 VSS.t1108 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X793 a_3822_2180.t0 a_3727_2165.t3 VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X794 a_2002_1924.t0 WWL[7].t7 a_2270_4887.t11 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X795 VSS.t499 a_5547_1698.t3 a_5452_1683.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X796 a_3727_2928.t0 WWL[3].t3 a_3995_4887.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X797 VDD.t1748 a_7847_2180.t4 a_7752_2165.t2 VDD.t1747 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X798 VSS.t452 a_2097_1216.t3 a_2002_1201.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X799 a_8452_n1770.t0 SA_OUT[14].t3 a_8360_n1371.t0 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X800 VDD.t5 SA_OUT[7].t3 a_4335_n1371.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X801 VSS.t1632 a_5547_n812.t3 a_5452_n827.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X802 a_3617_4445.t0 VSS.t718 a_3165_n953.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X803 VDD.t406 a_372_2180.t3 a_277_2165.t2 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X804 a_6133_n953.t20 WWL[13].t3 a_6122_452.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X805 a_7642_1216.t0 RWLB[10].t4 a_7190_n953.t36 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X806 VDD.t402 a_3493_n5850.t3 ADC6_OUT[1].t1 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X807 a_4302_3651.t2 WWL[0].t5 a_4570_4887.t23 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X808 a_947_2421.t2 a_852_2406.t3 VDD.t2112 VDD.t2111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X809 VSS.t996 a_1522_975.t3 a_1892_975.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X810 VDD.t1372 a_12963_n4483.t3 ADC14_OUT[0].t2 VDD.t1371 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X811 VSS.t2175 a_2672_n1053.t4 a_3042_n1053.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X812 a_7765_n953.t15 VSS.t717 a_7765_n512.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X813 a_6133_n953.t13 WWLD[2].t4 a_6122_4148.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X814 a_7283_n953.t20 WWL[6].t7 a_7272_2180.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X815 a_1427_1201.t0 WWL[10].t3 a_1695_4887.t8 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X816 a_4302_n45.t2 WWL[15].t3 a_4570_4887.t11 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X817 a_453_n2086.t1 WE.t8 a_383_n953.t12 VSS.t2381 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X818 a_8340_n953.t46 RWL[0].t4 a_8340_3666.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X819 a_8915_n953.t37 RWL[10].t6 a_8915_1216.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X820 VSS.t2321 a_6697_452.t3 a_7067_452.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X821 VSS.t2055 a_3247_n30.t3 a_3152_n45.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X822 a_947_n271.t1 a_852_n286.t3 VDD.t1324 VDD.t1323 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X823 a_8422_452.t0 a_8327_437.t3 VSS.t922 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X824 VDD.t1579 a_1522_1698.t3 a_1427_1683.t1 VDD.t1578 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X825 a_6040_n953.t46 RWL[12].t1 a_6040_693.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X826 a_8915_n1053.t1 a_8902_n1068.t3 VSS.t2466 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X827 a_865_n953.t1 RWL[0].t5 a_865_3666.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X828 a_3165_2180.t0 a_3152_2165.t5 VSS.t116 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X829 a_6727_n1770.t1 SA_OUT[11].t3 a_6635_n1371.t2 VSS.t1827 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X830 a_2015_4148.t1 a_2002_4133.t4 VSS.t229 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X831 VSS.t1623 a_4972_693.t3 a_4877_678.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X832 VDD.t2251 a_5547_693.t4 a_5452_678.t1 VDD.t2250 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X833 VSS.t1586 a_4397_3666.t3 a_4767_3666.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X834 a_5452_1924.t0 WWL[7].t8 a_5720_4887.t12 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X835 a_2311_n8583.t1 ADC5_OUT[3].t3 a_2381_n8071.t0 VSS.t1103 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X836 VDD.t804 a_2652_n2234.t2 a_2775_n2132.t1 VDD.t803 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X837 VDD.t1179 a_1522_n812.t3 a_1427_n827.t1 VDD.t1178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X838 a_3247_4148.t0 a_3152_4133.t3 VDD.t414 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X839 a_742_1939.t1 RWLB[7].t1 a_290_n953.t33 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X840 VSS.t1828 a_8422_452.t3 a_8792_452.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X841 VSS.t1043 a_4397_n512.t3 a_4302_n527.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X842 a_4890_n953.t12 VSS.t716 a_4890_4686.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X843 VSS.t450 a_4972_3666.t3 a_4877_3651.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X844 a_1317_3184.t1 RWLB[2].t2 a_865_n953.t48 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X845 VSS.t434 a_6122_1698.t3 a_6027_1683.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X846 VSS.t1561 a_5547_1216.t3 a_5452_1201.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X847 a_290_4445.t0 a_277_4430.t4 VSS.t2172 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X848 a_n2642_n5293.t1 VCLP.t18 a_n2677_n5092.t0 VSS.t180 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X849 a_4192_4445.t1 VSS.t715 a_3740_n953.t7 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X850 VSS.t776 a_6122_n812.t3 a_6027_n827.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X851 a_3740_n812.t1 a_3727_n827.t4 VSS.t2247 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X852 VSS.t1787 a_2672_1457.t4 a_3042_1457.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X853 a_13637_n5293.t1 VCLP.t19 a_13602_n5092.t0 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X854 a_6122_n812.t2 a_6027_n827.t3 VDD.t532 VDD.t531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X855 a_4397_2421.t2 a_4302_2406.t3 VDD.t1250 VDD.t1249 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 VSS.t1635 a_1522_4686.t3 a_1427_4671.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X857 a_5465_n953.t16 VSS.t714 a_5465_4445.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 a_8422_4445.t0 a_8327_4430.t3 VSS.t1571 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X859 a_4397_n271.t1 a_4302_n286.t3 VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X860 a_4302_n1068.t0 WWLD[7].t1 a_4570_4887.t25 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X861 a_8217_4686.t0 VSS.t713 a_7765_n953.t4 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X862 a_947_4445.t0 a_852_4430.t4 VSS.t64 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X863 a_1533_n953.t22 WWLD[7].t2 a_1522_n1053.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X864 a_6615_2180.t1 a_6602_2165.t4 VSS.t60 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X865 VSS.t1576 a_867_n4378.t4 a_867_n6849.t1 VSS.t1575 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X866 VDD.t1306 a_1522_1216.t3 a_1427_1201.t1 VDD.t1305 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 a_6027_n45.t0 WWL[15].t4 a_6295_4887.t24 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X868 a_7847_2180.t2 a_7752_2165.t3 VDD.t1023 VDD.t1022 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X869 a_2590_452.t0 a_2577_437.t4 VSS.t1974 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X870 a_6697_4148.t1 a_6602_4133.t3 VDD.t710 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X871 a_8902_3892.t0 WWLD[3].t5 a_9170_4887.t5 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X872 a_2108_n953.t23 WWL[8].t3 a_2097_1698.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X873 a_6027_1442.t2 WWL[9].t4 a_6295_4887.t20 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X874 a_5342_693.t1 RWLB[12].t1 a_4890_n953.t19 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X875 a_6812_n5293.t2 a_7039_n5850.t4 ADC9_OUT[1].t2 VSS.t429 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X876 VSS.t1519 a_2097_4445.t3 a_2002_4430.t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X877 a_4972_211.t2 a_4877_196.t4 VDD.t436 VDD.t435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X878 a_2590_n512.t1 a_2577_n527.t4 VSS.t2191 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X879 VDD.t1495 a_4972_3907.t3 a_4877_3892.t1 VDD.t1494 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X880 a_12963_n8583.t0 PRE_CLSA.t24 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X881 a_4972_n512.t2 a_4877_n527.t4 VDD.t1740 VDD.t1739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X882 a_7177_n1068.t0 WWLD[7].t3 a_7445_4887.t26 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X883 a_2108_n953.t17 WWLD[6].t5 a_2097_n812.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X884 a_277_2928.t0 WWL[3].t4 a_545_4887.t13 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X885 a_383_n953.t10 WWL[5].t2 a_372_2421.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X886 VSS.t1799 a_6122_1216.t3 a_6027_1201.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X887 a_7642_4445.t0 VSS.t712 a_7190_n953.t5 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X888 a_9178_n3770.t2 a_9405_n4483.t3 ADC11_OUT[0].t1 VSS.t1386 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X889 VSS.t1867 a_8997_3907.t3 a_9367_3907.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X890 a_3822_2662.t0 a_3727_2647.t3 VSS.t774 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X891 a_1120_4887.t8 WE.t9 a_1168_n2086.t1 VSS.t2382 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X892 VDD.t1624 a_6122_n1053.t3 a_6027_n1068.t1 VDD.t1623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X893 a_1427_4430.t2 WWLD[1].t3 a_1695_4887.t25 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X894 a_3247_4148.t1 a_3152_4133.t4 VSS.t480 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X895 a_3165_n953.t28 RWL[2].t5 a_3165_3184.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X896 a_6122_3184.t0 a_6027_3169.t3 VSS.t431 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X897 a_4397_2180.t0 a_4302_2165.t4 VSS.t476 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X898 VSS.t1915 a_6697_975.t4 a_7067_975.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X899 a_8915_n953.t5 VSS.t711 a_8915_4445.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X900 a_1533_n953.t20 WWL[13].t4 a_1522_452.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X901 VDD.t1515 a_5547_n30.t3 a_5452_n45.t1 VDD.t1514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X902 a_n2415_n5850.t1 ADC1_OUT[1].t3 VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X903 a_1533_n953.t23 WWL[9].t5 a_1522_1457.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X904 a_7765_975.t1 a_7752_960.t4 VSS.t2519 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X905 VDD.t2168 a_3822_n512.t4 a_3727_n527.t2 VDD.t2167 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X906 VSS.t1471 a_2097_452.t3 a_2467_452.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X907 a_3822_452.t1 a_3727_437.t3 VSS.t1453 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X908 a_5452_n1068.t0 WWLD[7].t4 a_5720_4887.t17 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X909 VDD.t1332 a_4397_3666.t4 a_4302_3651.t0 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X910 a_947_975.t1 a_852_960.t3 VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X911 a_1440_n953.t46 RWL[12].t2 a_1440_693.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X912 a_6040_4148.t1 a_6027_4133.t4 VSS.t2486 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X913 a_8997_2662.t1 a_8902_2647.t5 VDD.t1918 VDD.t1917 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X914 a_7190_2180.t1 a_7177_2165.t4 VSS.t2462 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X915 VDD.t1976 a_947_211.t4 a_852_196.t2 VDD.t1975 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X916 a_4972_n812.t0 a_4877_n827.t3 VSS.t240 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X917 VSS.t1595 a_5547_4445.t3 a_5452_4430.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X918 VSS.t465 a_8422_3666.t3 a_8792_3666.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X919 a_3995_4887.t15 WE.t10 a_4043_n2086.t0 VSS.t2383 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 a_2590_n953.t41 RWL[3].t2 a_2590_2943.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X921 VDD.t616 a_4972_n271.t3 a_4877_n286.t0 VDD.t615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X922 VSS.t969 a_8422_n512.t3 a_8327_n527.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X923 a_8902_3410.t0 WWL[1].t6 a_9170_4887.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X924 a_2108_n953.t9 WWL[10].t4 a_2097_1216.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X925 a_8422_n512.t2 a_8327_n527.t3 VDD.t1902 VDD.t1901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X926 a_2467_4148.t0 VSS.t710 a_2015_n953.t4 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X927 a_5342_3184.t1 RWLB[2].t3 a_4890_n953.t48 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X928 VSS.t1098 a_8997_n271.t3 a_9367_n271.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X929 VSS.t2356 a_9100_n2132.t2 a_9078_n2086.t1 VSS.t2355 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 a_2085_n1770.t0 PRE_VLSA.t10 VSS.t142 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X931 a_402_n1770.t0 a_383_n953.t27 a_360_n1770.t0 VSS.t803 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X932 VSS.t1777 a_2672_4686.t4 a_3042_4686.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X933 VDD.t942 a_4972_3425.t3 a_4877_3410.t2 VDD.t941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X934 VDD.t608 a_6122_1457.t3 a_6027_1442.t0 VDD.t607 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X935 a_1440_n953.t42 RWL[6].t1 a_1440_2180.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X936 a_7847_2180.t1 a_7752_2165.t4 VSS.t1670 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X937 a_6615_n953.t28 RWL[2].t6 a_6615_3184.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X938 a_8327_n1068.t0 WWLD[7].t5 a_8595_4887.t25 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X939 VSS.t1088 a_8997_3425.t3 a_9367_3425.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X940 a_6697_693.t2 a_6602_678.t3 VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X941 a_4675_n7216.t2 ADC7_OUT[2].t4 a_4745_n7203.t1 VSS.t1474 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X942 a_5145_4887.t19 PRE_SRAM.t11 VDD.t2031 VDD.t2030 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X943 a_7858_n953.t6 WWLD[3].t6 a_7847_3907.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X944 a_n52_n7216.t2 ADC3_OUT[2].t4 a_18_n7203.t2 VSS.t1083 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X945 a_3617_2421.t1 RWLB[5].t3 a_3165_n953.t48 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X946 a_5558_n953.t2 WWL[11].t9 a_5547_975.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X947 a_2270_4887.t9 WE.t11 a_2318_n2086.t0 VSS.t2384 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X948 VDD.t1273 a_1522_4445.t3 a_1427_4430.t0 VDD.t1272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X949 a_3617_n271.t0 VSS.t709 a_3165_n953.t11 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X950 VSS.t280 SAEN.t12 a_3266_n5293.t0 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X951 a_6027_4671.t0 WWLD[0].t4 a_6295_4887.t6 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X952 VSS.t1822 a_3247_3184.t3 a_3152_3169.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X953 a_2015_n953.t25 RWL[7].t1 a_2015_1939.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X954 VDD.t137 PRE_CLSA.t25 ADC14_OUT[2].t0 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X955 a_3247_n30.t1 a_3152_n45.t3 VSS.t1970 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X956 a_4408_n953.t4 WWLD[5].t8 a_4397_n512.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X957 a_1427_n45.t2 WWL[15].t5 a_1695_4887.t13 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X958 a_1129_n5850.t1 ADC4_OUT[1].t3 VDD.t1600 VDD.t827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X959 a_7067_n1053.t0 VSS.t708 a_6615_n953.t13 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X960 a_6133_n953.t1 WWL[8].t4 a_6122_1698.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X961 a_1502_n2234.t1 Din[2].t0 VDD.t1764 VDD.t1763 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X962 VSS.t1322 a_6122_4445.t3 a_6027_4430.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X963 a_5917_4148.t0 VSS.t707 a_5465_n953.t15 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X964 a_11984_n7203.t0 a_5743_n6391# a_11846_n7203.t2 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X965 VDD.t1630 a_8997_3907.t4 a_8902_3892.t1 VDD.t1629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X966 a_4972_n30.t0 a_4877_n45.t3 VSS.t1091 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X967 a_5145_4887.t24 WE.t12 a_5193_n2086.t1 VSS.t2385 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X968 a_2015_1698.t1 a_2002_1683.t4 VSS.t2467 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X969 a_n3792_n6503.t2 a_n3565_n7216.t4 ADC0_OUT[2].t2 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X970 a_6133_n953.t9 WWLD[6].t6 a_6122_n812.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X971 a_4890_n953.t27 RWL[4].t2 a_4890_2662.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X972 a_7858_n953.t9 WWLD[4].t6 a_7847_n271.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X973 a_1533_n953.t7 WWLD[0].t5 a_1522_4686.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X974 a_7272_4148.t1 a_7177_4133.t3 VSS.t1648 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X975 a_7190_n953.t0 RWL[2].t7 a_7190_3184.t1 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X976 a_3247_1698.t0 a_3152_1683.t3 VDD.t1540 VDD.t1539 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X977 a_742_n30.t1 RWLB[15].t3 a_290_n953.t36 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X978 a_4675_n7216.t0 PRE_CLSA.t26 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X979 a_7039_n8583.t1 ADC9_OUT[3].t3 a_7109_n8071.t2 VSS.t1939 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X980 VDD.t1505 a_5527_n2234.t2 a_5650_n2132.t1 VDD.t1504 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X981 a_2097_3666.t1 a_2002_3651.t3 VDD.t1546 VDD.t1545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X982 VSS.t2244 a_2672_2943.t3 a_2577_2928.t2 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X983 a_n1460_n6503.t1 VCLP.t20 a_n1495_n6849.t0 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X984 VDD.t141 PRE_CLSA.t27 ADC7_OUT[1].t0 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X985 a_290_2421.t0 a_277_2406.t4 VSS.t1063 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X986 a_n2207_n4470.t1 Iref0.t3 a_n2148_n4114.t1 VSS.t2219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X987 a_4377_n2234.t0 Din[7].t0 VDD.t1766 VDD.t1765 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X988 a_7858_n953.t0 WWL[1].t7 a_7847_3425.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X989 a_290_n271.t1 a_277_n286.t4 VSS.t2517 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X990 a_4192_2421.t1 RWLB[5].t4 a_3740_n953.t48 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X991 VSS.t282 SAEN.t13 a_11549_n8026.t0 VSS.t281 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X992 a_4192_n271.t0 VSS.t706 a_3740_n953.t20 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X993 VDD.t2183 a_13864_n5850.t3 ADC15_OUT[1].t2 VDD.t1036 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X994 VSS.t1662 a_1522_2662.t3 a_1427_2647.t0 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X995 a_5465_n953.t48 RWL[5].t6 a_5465_2421.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X996 a_8422_2421.t2 a_8327_2406.t3 VSS.t1278 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X997 a_1440_1457.t0 a_1427_1442.t4 VSS.t1202 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X998 a_12963_n5850.t2 ADC14_OUT[1].t4 a_13033_n5338.t2 VSS.t1484 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X999 a_2108_n953.t25 WWLD[1].t4 a_2097_4445.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1000 VSS.t2005 a_3822_3184.t3 a_3727_3169.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1001 VDD.t143 PRE_CLSA.t28 ADC3_OUT[0].t0 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1002 a_8217_2662.t0 RWLB[4].t0 a_7765_n953.t44 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1003 a_8422_n271.t0 a_8327_n286.t3 VSS.t1296 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1004 a_947_2421.t1 a_852_2406.t4 VSS.t2284 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1005 VDD.t714 a_8997_n271.t4 a_8902_n286.t2 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1006 VDD.t1867 a_6122_4686.t3 a_6027_4671.t2 VDD.t1866 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1007 a_947_n271.t0 a_852_n286.t4 VSS.t1569 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1008 VDD.t145 PRE_CLSA.t29 ADC2_OUT[1].t0 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1009 VDD.t638 a_8402_n2234.t2 a_8525_n2132.t1 VDD.t637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1010 a_6133_n953.t5 WWL[10].t5 a_6122_1216.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1011 a_2652_n2234.t0 Din[4].t0 VDD.t920 VDD.t919 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1012 a_8217_n1053.t0 VSS.t705 a_7765_n953.t6 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1013 a_6492_4148.t0 VSS.t704 a_6040_n953.t9 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1014 a_6602_3169.t0 WWL[2].t4 a_6870_4887.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1015 a_7858_n953.t23 WWL[13].t5 a_7847_452.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1016 a_8915_211.t0 a_8902_196.t3 VSS.t1058 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1017 VDD.t704 a_8997_3425.t4 a_8902_3410.t1 VDD.t703 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1018 a_7765_n953.t16 VSS.t703 a_7765_4148.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1019 a_1522_3907.t1 a_1427_3892.t3 VSS.t2109 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1020 VSS.t1326 a_2097_2421.t3 a_2002_2406.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1021 a_6697_1698.t2 a_6602_1683.t3 VDD.t1707 VDD.t1706 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1022 a_2015_1216.t1 a_2002_1201.t4 VSS.t799 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1023 a_2097_211.t1 a_2002_196.t3 VDD.t886 VDD.t885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1024 VDD.t1778 a_2672_3184.t3 a_2577_3169.t2 VDD.t1777 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1025 a_3822_2943.t1 a_3727_2928.t3 VSS.t1480 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1026 a_9170_4887.t22 PRE_SRAM.t12 VDD.t2033 VDD.t2032 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1027 a_3247_1216.t2 a_3152_1201.t3 VDD.t1709 VDD.t1708 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1028 a_9367_n812.t0 VSS.t702 a_8915_n953.t9 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1029 a_7642_2421.t0 RWLB[5].t5 a_7190_n953.t43 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1030 a_7272_975.t1 a_7177_960.t3 VDD.t1792 VDD.t1791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1031 a_2002_678.t2 WWL[12].t5 a_2270_4887.t7 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1032 VSS.t1650 a_1522_2180.t3 a_1892_2180.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1033 a_7765_n953.t32 RWL[12].t3 a_7765_693.t1 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1034 a_3152_n827.t0 WWLD[6].t7 a_3420_4887.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1035 a_1427_2406.t0 WWL[5].t3 a_1695_4887.t12 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1036 VDD.t59 a_7272_211.t4 a_7177_196.t2 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1037 a_7642_n271.t0 VSS.t701 a_7190_n953.t19 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1038 SA_OUT[13].t1 a_7785_n1371.t3 VDD.t1790 VDD.t1789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1039 a_7765_3907.t1 a_7752_3892.t5 VSS.t80 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1040 a_8915_n953.t34 RWL[5].t7 a_8915_2421.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1041 a_3247_1698.t1 a_3152_1683.t4 VSS.t1789 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1042 VSS.t1086 a_6697_693.t3 a_6602_678.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1043 a_1427_n286.t0 WWLD[4].t7 a_1695_4887.t16 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1044 a_5527_n2234.t0 Din[9].t0 VDD.t1857 VDD.t1856 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1045 VSS.t1328 a_4397_4148.t3 a_4302_4133.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1046 VSS.t1987 a_7272_3184.t3 a_7177_3169.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1047 a_6040_n953.t28 RWL[7].t2 a_6040_1939.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1048 a_4890_1939.t1 a_4877_1924.t5 VSS.t58 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1049 a_8433_n953.t7 WWLD[5].t9 a_8422_n512.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1050 a_8997_2943.t2 a_8902_2928.t5 VDD.t1302 VDD.t1301 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1051 a_7272_1939.t2 a_7177_1924.t3 VDD.t1169 VDD.t1168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1052 VSS.t1263 a_8422_211.t3 a_8327_196.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1053 a_958_n953.t3 WWLD[5].t10 a_947_n512.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1054 VSS.t2039 a_2097_1939.t3 a_2467_1939.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1055 VSS.t2097 a_8568_n2426.t4 a_12701_n5092.t1 VSS.t2095 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1056 VSS.t1335 a_5547_2421.t3 a_5452_2406.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1057 a_6040_1698.t1 a_6027_1683.t4 VSS.t2125 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1058 VSS.t1253 a_7847_2943.t3 a_7752_2928.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1059 a_11549_n5293.t1 VCLP.t21 a_11514_n5092.t0 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1060 a_4675_n4483.t0 ADC7_OUT[0].t3 a_4745_n4470.t0 VSS.t1262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1061 a_2002_n527.t2 WWLD[5].t11 a_2270_4887.t4 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1062 a_2672_1457.t1 a_2577_1442.t3 VSS.t1962 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1063 a_n52_n4483.t1 ADC3_OUT[0].t3 a_18_n4470.t2 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1064 a_1522_3425.t1 a_1427_3410.t3 VSS.t2037 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1065 a_6697_1216.t1 a_6602_1201.t3 VDD.t1521 VDD.t1520 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1066 VDD.t375 a_8997_452.t4 a_8902_437.t0 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1067 VSS.t985 a_6693_n2422.t4 a_9143_n6849.t0 VSS.t984 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1068 VSS.t918 a_2672_2662.t4 a_3042_2662.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1069 a_2467_1698.t1 RWLB[8].t5 a_2015_n953.t31 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1070 a_2590_n1053.t1 a_2577_n1068.t4 VSS.t2336 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1071 a_1317_3666.t0 RWLB[0].t2 a_865_n953.t26 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1072 a_1440_4686.t1 a_1427_4671.t4 VSS.t778 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1073 a_7067_211.t1 RWLB[14].t3 a_6615_n953.t43 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1074 VDD.t2035 PRE_SRAM.t13 a_6708_n953.t23 VDD.t2034 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1075 a_11776_n8583.t2 ADC13_OUT[3].t3 VDD.t848 VDD.t847 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1076 a_6615_n953.t42 EN.t0 a_6693_n2422.t2 VSS.t2041 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1077 a_7765_3425.t1 a_7752_3410.t5 VSS.t2162 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1078 a_3247_1216.t0 a_3152_1201.t4 VSS.t999 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1079 a_8997_975.t1 a_8902_960.t3 VDD.t422 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1080 a_3727_678.t2 WWL[12].t6 a_3995_4887.t10 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1081 SA_OUT[15].t1 a_8935_n1371.t3 VDD.t620 VDD.t619 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1082 a_6133_n953.t16 WWLD[1].t5 a_6122_4445.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1083 VDD.t1422 a_1522_2421.t3 a_1427_2406.t2 VDD.t1421 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1084 a_9405_n5850.t0 PRE_CLSA.t30 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1085 a_11984_n4470.t0 VCLP.t22 a_11846_n4470.t2 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1086 a_6027_2647.t2 WWL[4].t4 a_6295_4887.t21 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1087 VSS.t1682 a_5547_1939.t3 a_5917_1939.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1088 a_372_1457.t2 a_277_1442.t3 VDD.t564 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1089 a_8792_211.t1 RWLB[14].t4 a_8340_n953.t36 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1090 VDD.t420 a_n1233_n8583.t3 ADC2_OUT[3].t1 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1091 a_n3792_n3770.t2 a_n3565_n4483.t3 ADC0_OUT[0].t2 VSS.t427 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1092 a_2015_4445.t1 a_2002_4430.t4 VSS.t1092 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1093 a_1892_1457.t1 RWLB[9].t1 a_1440_n953.t31 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1094 a_7272_693.t1 a_7177_678.t3 VSS.t2181 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1095 a_290_452.t0 a_277_437.t4 VSS.t443 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1096 a_7835_n1770.t0 PRE_VLSA.t11 VSS.t146 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1097 a_5452_n527.t2 WWLD[5].t12 a_5720_4887.t4 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1098 a_3247_4445.t1 a_3152_4430.t3 VDD.t1817 VDD.t1816 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1099 a_2590_n953.t13 VSS.t700 a_2590_3907.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1100 a_8997_3907.t0 a_8902_3892.t4 VSS.t1291 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1101 VSS.t1476 a_6122_2421.t3 a_6027_2406.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1102 a_6040_1216.t0 a_6027_1201.t4 VSS.t1610 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 a_742_n512.t0 VSS.t699 a_290_n953.t10 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1104 a_n1460_n3770.t1 VCLP.t23 a_n1495_n4116.t0 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1105 VDD.t686 a_3822_4148.t4 a_3727_4133.t1 VDD.t685 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1106 VDD.t1312 a_6697_3184.t3 a_6602_3169.t1 VDD.t1311 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1107 a_5917_1698.t1 RWLB[8].t6 a_5465_n953.t34 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1108 a_3042_975.t0 RWLB[11].t4 a_2590_n953.t43 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1109 VSS.t49 a_6697_2180.t4 a_7067_2180.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1110 a_3165_n953.t47 RWL[14].t3 a_3165_211.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1111 a_7177_n827.t0 WWLD[6].t8 a_7445_4887.t8 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1112 a_2467_1216.t0 RWLB[10].t5 a_2015_n953.t37 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1113 a_2672_975.t2 a_2577_960.t3 VDD.t1650 VDD.t1649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1114 a_3740_n1053.t1 a_3727_n1068.t4 VSS.t2465 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1115 a_1533_n953.t24 WWL[4].t5 a_1522_2662.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1116 a_4315_452.t1 a_4302_437.t4 VSS.t1314 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1117 VSS.t2023 a_2097_211.t3 a_2002_196.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1118 VDD.t1936 a_2672_211.t4 a_2577_196.t1 VDD.t1935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1119 a_1552_n1770.t1 SA_OUT[2].t3 a_1460_n1371.t2 VSS.t2493 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1120 a_7272_1698.t2 a_7177_1683.t3 VSS.t1819 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1121 VDD.t2261 a_11776_n4483.t4 ADC13_OUT[0].t1 VDD.t2260 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1122 VSS.t1896 a_8422_4148.t3 a_8327_4133.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1123 a_3165_n953.t29 RWL[0].t6 a_3165_3666.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1124 a_6122_3666.t0 a_6027_3651.t3 VSS.t1584 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1125 VDD.t1646 a_2311_n7216.t3 ADC5_OUT[2].t2 VDD.t797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1126 VDD.t1483 a_7272_2943.t3 a_7177_2928.t2 VDD.t1482 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1127 VDD.t1794 a_2097_1939.t4 a_2002_1924.t1 VDD.t1793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1128 a_4890_n953.t24 RWL[14].t4 a_4890_211.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1129 VSS.t283 SAEN.t14 a_13637_n5293.t0 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1130 a_7765_n953.t46 EN.t1 a_7843_n2422.t3 VSS.t2042 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1131 a_8217_2943.t1 RWLB[3].t0 a_7765_n953.t43 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1132 a_3042_1939.t1 RWLB[7].t2 a_2590_n953.t33 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1133 VSS.t1541 a_6122_1939.t3 a_6492_1939.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1134 a_n1233_n4483.t2 ADC2_OUT[0].t4 VDD.t544 VDD.t543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1135 a_2108_n953.t6 WWL[5].t4 a_2097_2421.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1136 a_2590_n953.t12 VSS.t698 a_2590_n271.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1137 a_2672_4686.t2 a_2577_4671.t3 VSS.t1967 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1138 a_947_3184.t1 a_852_3169.t3 VDD.t588 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1139 a_8422_211.t1 a_8327_196.t3 VDD.t1683 VDD.t1682 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1140 a_6697_4445.t1 a_6602_4430.t3 VDD.t722 VDD.t721 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1141 VDD.t1463 a_6122_n30.t4 a_6027_n45.t2 VDD.t1462 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1142 VSS.t1135 a_372_2943.t3 a_742_2943.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1143 VDD.t1491 a_6122_2662.t3 a_6027_2647.t0 VDD.t1490 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1144 a_3740_n953.t26 RWL[11].t1 a_3740_975.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1145 a_8429_n7203.t0 a_5743_n6391# a_8291_n7203.t2 VSS.t225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1146 a_4983_n953.t24 WWL[15].t6 a_4972_n30.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1147 a_2590_n953.t21 RWL[1].t2 a_2590_3425.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1148 a_8997_3425.t1 a_8902_3410.t4 VSS.t1431 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1149 a_10589_n4483.t0 PRE_CLSA.t31 VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1150 VSS.t1451 a_3822_452.t3 a_3727_437.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1151 a_5342_3666.t0 RWLB[0].t3 a_4890_n953.t28 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1152 a_6492_1698.t1 RWLB[8].t7 a_6040_n953.t34 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1153 a_5917_1216.t0 RWLB[10].t6 a_5465_n953.t40 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1154 VDD.t1378 a_4397_452.t4 a_4302_437.t2 VDD.t1377 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1155 a_n1025_n8071.t1 Iref3.t3 a_n966_n8026.t1 VSS.t1983 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1156 VSS.t285 SAEN.t15 a_5630_n8026.t0 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1157 VSS.t1963 a_947_n1053.t3 a_1317_n1053.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1158 a_4408_n953.t17 WWLD[2].t5 a_4397_4148.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1159 a_5558_n953.t25 WWL[6].t8 a_5547_2180.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 a_3247_4445.t2 a_3152_4430.t4 VSS.t2070 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1161 VSS.t1890 a_2672_3907.t3 a_2577_3892.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1162 a_6615_n953.t29 RWL[0].t7 a_6615_3666.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1163 a_7765_n953.t42 RWL[8].t5 a_7765_1698.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1164 a_2467_211.t1 RWLB[14].t5 a_2015_n953.t38 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1165 a_372_4686.t1 a_277_4671.t3 VDD.t1275 VDD.t1274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1166 VDD.t1424 a_5547_1939.t4 a_5452_1924.t1 VDD.t1423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1167 VSS.t493 a_5547_452.t3 a_5917_452.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1168 VSS.t287 SAEN.t16 a_7994_n8026.t0 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1169 a_7272_1216.t2 a_7177_1201.t3 VSS.t1897 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1170 a_4397_975.t1 a_4302_960.t3 VDD.t1863 VDD.t1862 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1171 a_7765_n953.t17 VSS.t697 a_7765_n812.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1172 a_1892_4686.t0 VSS.t696 a_1440_n953.t16 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1173 a_7067_1457.t0 RWLB[9].t2 a_6615_n953.t36 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1174 a_2381_n7203.t0 SAEN.t17 a_2578_n6847.t0 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1175 a_1522_4148.t1 a_1427_4133.t3 VDD.t1599 VDD.t1598 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1176 a_4397_3184.t2 a_4302_3169.t3 VDD.t960 VDD.t959 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1177 a_2672_2180.t1 a_2577_2165.t3 VDD.t1616 VDD.t1615 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1178 a_852_1442.t2 WWL[9].t6 a_1120_4887.t16 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1179 a_6040_4445.t1 a_6027_4430.t4 VSS.t1324 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1180 a_3266_n5293.t1 a_3493_n5850.t4 ADC6_OUT[1].t2 VSS.t461 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1181 VSS.t261 a_3247_3666.t5 a_3152_3651.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1182 VSS.t407 a_4397_1698.t5 a_4302_1683.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1183 a_2672_693.t1 a_2577_678.t3 VSS.t150 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1184 a_5465_n30.t1 a_5452_n45.t4 VSS.t1972 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1185 a_4983_n953.t16 WWL[7].t9 a_4972_1939.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1186 VSS.t288 SAEN.t18 a_6812_n5293.t0 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1187 VDD.t151 PRE_CLSA.t32 ADC5_OUT[2].t0 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1188 a_11776_n8583.t0 PRE_CLSA.t33 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1189 a_2467_4445.t0 VSS.t695 a_2015_n953.t5 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1190 VSS.t236 a_4397_n812.t5 a_4302_n827.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1191 a_372_1939.t0 a_277_1924.t3 VSS.t456 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1192 VSS.t1189 a_947_1457.t3 a_1317_1457.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1193 VSS.t1694 a_1050_n2132.t2 a_1028_n2086.t1 VSS.t1693 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1194 a_4192_452.t0 RWLB[13].t3 a_3740_n953.t25 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1195 VSS.t1182 a_2672_n271.t3 a_2577_n286.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1196 a_6492_1216.t0 RWLB[10].t7 a_6040_n953.t40 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1197 a_5558_n953.t22 WWL[15].t7 a_5547_n30.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1198 VSS.t1023 a_n2677_n4378.t5 a_n2677_n4116.t1 VSS.t1019 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1199 a_7190_n953.t1 RWL[0].t8 a_7190_3666.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1200 VSS.t1555 a_2672_3425.t3 a_2577_3410.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1201 a_7765_n953.t38 RWL[10].t7 a_7765_1216.t1 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1202 VSS.t1505 a_4397_n30.t3 a_4767_n30.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1203 VDD.t1536 a_n52_n4483.t4 ADC3_OUT[0].t1 VDD.t1535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1204 a_383_n953.t1 WWL[2].t5 a_372_3184.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1205 a_1440_2662.t0 a_1427_2647.t4 VSS.t1666 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1206 a_3727_3892.t0 WWLD[3].t7 a_3995_4887.t9 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1207 a_865_975.t1 a_852_960.t4 VSS.t849 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1208 VDD.t155 PRE_CLSA.t34 ADC6_OUT[0].t0 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1209 a_6027_2928.t0 WWL[3].t5 a_6295_4887.t18 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1210 a_4302_1924.t0 WWL[7].t10 a_4570_4887.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1211 SA_OUT[13].t0 PRE_VLSA.t12 VDD.t1149 VDD.t1148 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1212 a_6133_n953.t3 WWL[5].t5 a_6122_2421.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1213 a_5630_n5293.t1 VCLP.t24 a_5595_n5092.t0 VSS.t186 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1214 a_9367_975.t1 RWLB[11].t5 a_8915_n953.t20 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1215 a_3822_211.t2 a_3727_196.t3 VDD.t818 VDD.t817 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1216 a_2084_n6503.t1 VCLP.t25 a_2049_n6849.t0 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1217 VSS.t2421 a_3822_3666.t4 a_3727_3651.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1218 VSS.t2417 a_4397_1216.t5 a_4302_1201.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1219 VDD.t1002 a_2097_n30.t3 a_2002_n45.t2 VDD.t1001 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1220 a_5917_4445.t0 VSS.t694 a_5465_n953.t14 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1221 a_2015_2421.t0 a_2002_2406.t4 VSS.t488 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1222 VDD.t1724 a_947_n1053.t4 a_852_n1068.t1 VDD.t1723 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1223 VSS.t1130 a_2672_693.t3 a_3042_693.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1224 a_2015_n271.t1 a_2002_n286.t4 VSS.t2149 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1225 a_2590_n812.t1 a_2577_n827.t4 VSS.t1345 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1226 VSS.t2358 a_7847_3907.t5 a_7752_3892.t2 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1227 a_4972_n812.t1 a_4877_n827.t4 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1228 a_6602_3651.t2 WWL[0].t6 a_6870_4887.t26 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1229 a_3247_2421.t2 a_3152_2406.t3 VDD.t1603 VDD.t1602 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1230 VSS.t1643 a_2200_n2132.t2 a_2178_n2086.t1 VSS.t1642 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 VSS.t2409 a_4972_n1053.t4 a_5342_n1053.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1232 a_7272_4445.t1 a_7177_4430.t3 VSS.t1861 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1233 a_8433_n953.t23 WWLD[2].t6 a_8422_4148.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1234 a_3247_n271.t1 a_3152_n286.t3 VDD.t996 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1235 a_5857_n8583.t1 ADC8_OUT[3].t3 VDD.t790 VDD.t789 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1236 VDD.t950 a_3822_1698.t4 a_3727_1683.t2 VDD.t949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1237 VSS.t2364 a_8997_n1053.t5 a_8902_n1068.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1238 a_7067_4686.t0 VSS.t693 a_6615_n953.t9 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1239 a_958_n953.t14 WWLD[2].t7 a_947_4148.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1240 VDD.t1968 a_2672_3666.t3 a_2577_3651.t1 VDD.t1967 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1241 VDD.t157 PRE_CLSA.t35 ADC4_OUT[3].t0 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1242 a_1427_n1068.t1 WWLD[7].t6 a_1695_4887.t22 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1243 a_852_4671.t0 WWLD[0].t6 a_1120_4887.t24 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1244 a_4315_4148.t1 a_4302_4133.t4 VSS.t1817 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1245 a_5465_2180.t0 a_5452_2165.t5 VSS.t1821 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1246 VDD.t1263 a_4675_n7216.t3 ADC7_OUT[2].t1 VDD.t1084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1247 a_5547_452.t0 a_5452_437.t3 VDD.t787 VDD.t786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1248 VDD.t1920 a_3822_n812.t4 a_3727_n827.t1 VDD.t1919 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1249 VSS.t2511 a_6697_n512.t4 a_6602_n527.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1250 a_5547_4148.t0 a_5452_4133.t3 VDD.t580 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 a_3727_3410.t0 WWL[1].t8 a_3995_4887.t2 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1252 a_4877_1442.t0 WWL[9].t7 a_5145_4887.t13 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1253 VSS.t2334 a_7272_3666.t4 a_7177_3651.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1254 VSS.t2170 a_8422_1698.t4 a_8327_1683.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1255 a_n2415_n5850.t2 ADC1_OUT[1].t4 a_n2345_n5338.t1 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1256 a_8429_n4470.t0 VCLP.t26 a_8291_n4470.t1 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1257 a_3617_3184.t1 RWLB[2].t4 a_3165_n953.t45 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1258 VSS.t1878 a_947_4686.t3 a_1317_4686.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1259 VDD.t820 a_947_1457.t4 a_852_1442.t0 VDD.t819 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1260 a_4972_n1053.t1 a_4877_n1068.t3 VDD.t2178 VDD.t2177 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1261 a_4397_n1053.t0 a_4302_n1068.t4 VSS.t2443 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1262 SA_OUT[15].t2 PRE_VLSA.t13 VDD.t1147 VDD.t1146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1263 VSS.t2246 a_7847_n271.t5 a_7752_n286.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1264 VSS.t1497 a_5632_n6430# a_12736_n6503.t0 VSS.t273 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1265 VSS.t2214 a_8422_n812.t4 a_8327_n827.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1266 a_6492_4445.t0 VSS.t692 a_6040_n953.t5 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1267 a_8422_n812.t1 a_8327_n827.t3 VDD.t1175 VDD.t1174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1268 a_2672_2662.t1 a_2577_2647.t3 VSS.t1832 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1269 a_6697_2421.t2 a_6602_2406.t3 VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1270 VSS.t2216 a_4972_1457.t4 a_5342_1457.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1271 a_3493_n8583.t1 ADC6_OUT[3].t3 a_3563_n8071.t2 VSS.t1424 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1272 a_12963_n5850.t0 PRE_CLSA.t36 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1273 a_2097_4148.t0 a_2002_4133.t5 VSS.t114 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1274 a_7765_n953.t13 VSS.t691 a_7765_4445.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1275 a_6697_n271.t0 a_6602_n286.t3 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1276 VSS.t2455 a_2049_n4378.t4 a_2049_n5092.t1 VSS.t2453 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1277 VDD.t1750 a_5857_n4483.t4 ADC8_OUT[0].t2 VDD.t1749 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1278 VSS.t2310 a_7847_3425.t5 a_7752_3410.t2 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1279 VSS.t2307 a_8997_1457.t5 a_8902_1442.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1280 a_1533_n953.t13 WWL[15].t8 a_1522_n30.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1281 a_n3565_n7216.t1 ADC0_OUT[2].t3 VDD.t365 VDD.t364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1282 a_5452_678.t2 WWL[12].t7 a_5720_4887.t8 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1283 a_3833_n953.t20 WWLD[7].t7 a_3822_n1053.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1284 a_8915_2180.t0 a_8902_2165.t3 VSS.t1859 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1285 VSS.t290 SAEN.t19 a_10362_n8026.t0 VSS.t289 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1286 VDD.t1477 a_3822_1216.t4 a_3727_1201.t1 VDD.t1476 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1287 a_2381_n4470.t0 SAEN.t20 a_2578_n4114.t0 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1288 a_3247_2421.t1 a_3152_2406.t4 VSS.t1848 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1289 a_7177_196.t0 WWL[14].t10 a_7445_4887.t19 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1290 VDD.t1728 a_8221_n4483.t4 ADC10_OUT[0].t1 VDD.t1727 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1291 a_927_n2234.t0 Din[1].t1 VSS.t2524 VSS.t2523 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1292 a_7272_n1053.t1 a_7177_n1068.t3 VSS.t1903 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1293 a_8327_1442.t2 WWL[9].t8 a_8595_4887.t16 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1294 a_8997_693.t1 a_8902_678.t3 VSS.t1120 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1295 a_3042_n1053.t1 VSS.t690 a_2590_n953.t18 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1296 a_4408_n953.t2 WWL[8].t5 a_4397_1698.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1297 a_3247_n271.t2 a_3152_n286.t4 VSS.t1360 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1298 VSS.t2429 a_4397_4445.t5 a_4302_4430.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1299 a_372_2662.t1 a_277_2647.t3 VDD.t353 VDD.t352 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1300 a_4972_n30.t1 a_4877_n45.t4 VDD.t912 VDD.t911 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1301 a_4745_n7203.t0 SAEN.t21 a_4942_n6847.t0 VSS.t275 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1302 a_277_3892.t0 WWLD[3].t8 a_545_4887.t6 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1303 a_290_3184.t0 a_277_3169.t4 VSS.t1696 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1304 a_4890_n512.t1 a_4877_n527.t5 VSS.t811 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1305 VDD.t2006 a_7272_3907.t3 a_7177_3892.t2 VDD.t2005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1306 a_1892_2662.t1 RWLB[4].t1 a_1440_n953.t35 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1307 a_7272_n512.t1 a_7177_n527.t3 VDD.t1906 VDD.t1905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1308 a_4192_3184.t0 RWLB[2].t5 a_3740_n953.t4 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1309 VSS.t2331 a_8422_1216.t4 a_8327_1201.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1310 a_4767_975.t0 RWLB[11].t6 a_4315_n953.t43 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1311 VDD.t1762 a_4972_975.t3 a_4877_960.t1 VDD.t1761 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1312 a_4408_n953.t12 WWLD[6].t9 a_4397_n812.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1313 VDD.t1693 a_8422_n1053.t3 a_8327_n1068.t1 VDD.t1692 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1314 a_5547_4148.t1 a_5452_4133.t4 VSS.t933 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1315 a_6040_2421.t0 a_6027_2406.t4 VSS.t1050 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1316 a_6697_2180.t0 a_6602_2165.t5 VSS.t65 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1317 a_1522_1698.t1 a_1427_1683.t3 VDD.t946 VDD.t945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1318 VSS.t1268 a_8997_975.t3 a_9367_975.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1319 a_7109_n7203.t0 a_5632_n6430# a_7306_n6847.t0 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1320 a_5465_n953.t27 RWL[2].t8 a_5465_3184.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1321 a_8422_3184.t0 a_8327_3169.t4 VSS.t404 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1322 a_6040_n271.t1 a_6027_n286.t4 VSS.t1032 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1323 a_1129_n5850.t2 ADC4_OUT[1].t4 a_1199_n5338.t2 VSS.t1638 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1324 VDD.t2092 a_1502_n2234.t3 a_1625_n2132.t1 VDD.t2091 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1325 a_6122_n1053.t1 a_6027_n1068.t3 VDD.t1638 VDD.t1637 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1326 a_5547_n1053.t0 a_5452_n1068.t3 VSS.t766 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1327 VSS.t2320 a_372_3907.t4 a_742_3907.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1328 a_1317_n1053.t0 VSS.t689 a_865_n953.t17 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1329 a_947_3184.t2 a_852_3169.t4 VSS.t940 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1330 a_958_n953.t21 WWL[13].t6 a_947_452.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1331 a_3995_4887.t5 PRE_SRAM.t14 VDD.t2037 VDD.t2036 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1332 a_3833_n953.t21 WWL[9].t9 a_3822_1457.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1333 a_2467_2421.t1 RWLB[5].t6 a_2015_n953.t43 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1334 a_2467_n271.t0 VSS.t688 a_2015_n953.t16 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1335 VSS.t1931 a_7847_n512.t3 a_8217_n512.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1336 VDD.t1703 a_6697_3666.t3 a_6602_3651.t0 VDD.t1702 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1337 a_4877_4671.t2 WWLD[0].t7 a_5145_4887.t18 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1338 a_2108_n953.t22 WWL[15].t9 a_2097_n30.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1339 a_8340_4148.t1 a_8327_4133.t4 VSS.t1227 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1340 VSS.t2508 a_2097_3184.t5 a_2002_3169.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1341 a_372_975.t1 a_277_960.t3 VDD.t844 VDD.t843 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1342 a_2519_n8071.t0 VCLP.t27 a_2381_n8071.t2 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1343 a_865_n953.t42 RWL[12].t4 a_865_693.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1344 a_8433_n953.t11 WWL[12].t8 a_8422_693.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1345 a_3258_n953.t2 WWLD[5].t13 a_3247_n512.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1346 a_865_4148.t1 a_852_4133.t5 VSS.t1993 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1347 a_1440_2943.t1 a_1427_2928.t4 VSS.t1479 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1348 VDD.t1454 a_372_211.t4 a_277_196.t2 VDD.t1453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1349 VSS.t1607 a_947_n30.t3 a_1317_n30.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1350 VDD.t2158 a_7272_n271.t3 a_7177_n286.t1 VDD.t2157 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1351 VDD.t736 a_947_4686.t4 a_852_4671.t1 VDD.t735 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1352 a_4890_n953.t17 RWL[3].t3 a_4890_2943.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1353 a_2084_n3770.t1 VCLP.t28 a_2049_n4116.t0 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1354 SA_OUT[8].t1 a_4910_n1371.t3 a_5153_n1770.t1 VSS.t1458 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1355 SA_OUT[1].t2 a_885_n1371.t3 VDD.t1699 VDD.t1698 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1356 a_8422_n1053.t1 a_8327_n1068.t3 VSS.t963 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1357 a_4408_n953.t5 WWL[10].t6 a_4397_1216.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1358 a_8997_n1053.t2 a_8902_n1068.t4 VDD.t2229 VDD.t2228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1359 a_4767_4148.t0 VSS.t687 a_4315_n953.t14 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1360 a_7642_3184.t1 RWLB[2].t6 a_7190_n953.t45 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1361 a_5857_n8583.t0 PRE_CLSA.t37 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1362 a_277_3410.t2 WWL[1].t9 a_545_4887.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1363 VDD.t1063 a_8422_1457.t3 a_8327_1442.t0 VDD.t1062 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1364 VSS.t1118 a_8997_693.t3 a_9367_693.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1365 a_8340_n953.t35 EN.t2 a_8568_n2426.t2 VSS.t2043 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1366 VSS.t2491 a_4972_4686.t4 a_5342_4686.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1367 VDD.t412 a_7272_3425.t3 a_7177_3410.t2 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1368 a_1427_3169.t0 WWL[2].t6 a_1695_4887.t3 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1369 a_4448_n6503.t2 VCLP.t29 a_4413_n6849.t0 VSS.t164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1370 a_5193_n2086.t0 a_4952_n2234.t3 VSS.t1248 VSS.t1247 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1371 a_8915_n953.t28 RWL[2].t9 a_8915_3184.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1372 a_3740_n953.t44 RWL[6].t2 a_3740_2180.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1373 VSS.t2489 a_372_n271.t4 a_742_n271.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1374 a_13637_n5293.t2 a_13864_n5850.t4 ADC15_OUT[1].t1 VSS.t1236 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1375 VDD.t163 PRE_CLSA.t38 ADC10_OUT[0].t0 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1376 VSS.t2285 a_8997_4686.t5 a_8902_4671.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1377 a_10362_n5293.t1 VCLP.t30 a_10327_n5092.t0 VSS.t190 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1378 a_7445_4887.t21 PRE_SRAM.t15 VDD.t2039 VDD.t2038 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1379 a_947_3666.t0 a_852_3651.t3 VDD.t1025 VDD.t1024 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 VSS.t798 a_1522_2943.t4 a_1427_2928.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1381 a_1522_1216.t2 a_1427_1201.t3 VDD.t1281 VDD.t1280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1382 a_5917_2421.t0 RWLB[5].t7 a_5465_n953.t44 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1383 a_7858_n953.t1 WWL[11].t10 a_7847_975.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1384 a_n2642_n8026.t2 a_n2415_n8583.t3 ADC1_OUT[3].t2 VSS.t1416 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1385 VSS.t2272 a_372_3425.t4 a_742_3425.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1386 a_852_196.t0 WWL[14].t11 a_1120_4887.t11 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1387 a_6615_n953.t48 RWL[14].t5 a_6615_211.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1388 SA_OUT[5].t1 a_3185_n1371.t3 a_3428_n1770.t1 VSS.t2420 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1389 a_9008_n953.t26 WWLD[7].t8 a_8997_n1053.t1 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1390 VDD.t674 a_3822_4445.t4 a_3727_4430.t1 VDD.t673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1391 a_5917_n271.t0 VSS.t686 a_5465_n953.t6 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1392 VSS.t293 SAEN.t22 a_902_n8026.t0 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1393 SA_OUT[6].t0 a_3760_n1371.t3 VDD.t1320 VDD.t1319 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1394 a_8327_4671.t0 WWLD[0].t8 a_8595_4887.t20 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1395 VSS.t67 a_5547_211.t3 a_5452_196.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1396 VSS.t475 a_5547_3184.t5 a_5452_3169.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1397 a_4315_n953.t25 RWL[7].t3 a_4315_1939.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1398 a_4397_211.t1 a_4302_196.t3 VSS.t1785 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1399 a_8068_n2086.t1 a_7827_n2234.t3 VSS.t406 VSS.t405 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1400 a_6708_n953.t2 WWLD[5].t14 a_6697_n512.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1401 a_7272_2421.t1 a_7177_2406.t4 VSS.t2378 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1402 a_2097_1939.t1 a_2002_1924.t3 VDD.t1461 VDD.t1460 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1403 a_2577_196.t2 WWL[14].t12 a_2845_4887.t17 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1404 a_10589_n8583.t1 ADC12_OUT[3].t3 VDD.t1318 VDD.t1317 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1405 a_8433_n953.t5 WWL[8].t6 a_8422_1698.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1406 a_7272_n271.t0 a_7177_n286.t4 VSS.t2351 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1407 VSS.t1211 a_5543_n2422.t5 a_6777_n4116.t1 VSS.t1207 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1408 VSS.t796 a_8422_4445.t4 a_8327_4430.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1409 a_7067_2662.t1 RWLB[4].t2 a_6615_n953.t40 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1410 a_852_2647.t2 WWL[4].t6 a_1120_4887.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1411 a_3165_693.t1 a_3152_678.t4 VSS.t790 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1412 a_958_n953.t1 WWL[8].t7 a_947_1698.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1413 a_2660_n1770.t0 PRE_VLSA.t14 VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1414 a_4315_1698.t1 a_4302_1683.t4 VSS.t2252 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1415 VDD.t902 a_8997_975.t4 a_8902_960.t1 VDD.t901 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1416 VSS.t295 SAEN.t23 a_12736_n3770.t0 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1417 VDD.t165 PRE_CLSA.t39 ADC15_OUT[0].t0 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1418 a_8433_n953.t17 WWLD[6].t10 a_8422_n812.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1419 VSS.t974 a_947_1939.t5 a_852_1924.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1420 a_2311_n7216.t1 ADC5_OUT[2].t3 VDD.t1645 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1421 SA_OUT[10].t0 a_6060_n1371.t3 a_6303_n1770.t1 VSS.t869 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1422 SA_OUT[3].t2 a_2035_n1371.t3 VDD.t327 VDD.t326 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1423 a_3042_n512.t0 VSS.t685 a_2590_n953.t10 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1424 a_958_n953.t10 WWLD[6].t11 a_947_n812.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1425 a_3833_n953.t7 WWLD[0].t9 a_3822_4686.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1426 a_4397_3666.t1 a_4302_3651.t3 VDD.t1279 VDD.t1278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1427 a_5547_1698.t0 a_5452_1683.t3 VDD.t393 VDD.t392 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1428 a_8340_n953.t37 RWL[13].t2 a_8340_452.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1429 a_6343_n2086.t1 a_6102_n2234.t2 VSS.t864 VSS.t863 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1430 a_9008_n953.t11 WWL[9].t10 a_8997_1457.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1431 a_372_693.t2 a_277_678.t3 VSS.t2330 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1432 a_4890_693.t0 a_4877_678.t3 VSS.t1621 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1433 VDD.t1489 a_1522_3184.t3 a_1427_3169.t1 VDD.t1488 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1434 a_2672_2943.t1 a_2577_2928.t4 VSS.t2251 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1435 VSS.t1753 a_947_2662.t3 a_1317_2662.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1436 VDD.t1701 a_7847_n512.t4 a_7752_n527.t2 VDD.t1700 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1437 VSS.t464 a_7272_452.t3 a_7177_437.t0 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1438 a_6492_2421.t1 RWLB[5].t8 a_6040_n953.t43 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 a_2108_n953.t11 WWL[12].t9 a_2097_693.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1440 VDD.t2138 a_372_n512.t3 a_277_n527.t2 VDD.t2137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1441 VSS.t396 a_7950_n2132.t2 a_7928_n2086.t1 VSS.t395 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1442 a_2002_n827.t0 WWLD[6].t12 a_2270_4887.t13 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1443 a_6492_n271.t0 VSS.t684 a_6040_n953.t2 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1444 a_8429_n4470.t1 Iref0.t4 a_8488_n4114.t1 VSS.t2220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1445 a_7765_n953.t36 RWL[5].t8 a_7765_2421.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 a_5917_211.t1 RWLB[14].t6 a_5465_n953.t41 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1447 SA_OUT[7].t1 a_4335_n1371.t3 a_4578_n1770.t0 VSS.t1461 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1448 a_2097_1698.t0 a_2002_1683.t5 VSS.t2468 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1449 a_3740_1457.t0 a_3727_1442.t4 VSS.t2137 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1450 a_14072_n8071.t1 Iref3.t4 a_14131_n8026.t1 VSS.t1984 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1451 VDD.t1568 a_10589_n4483.t4 ADC12_OUT[0].t2 VDD.t1567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1452 a_4408_n953.t18 WWLD[1].t6 a_4397_4445.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1453 VSS.t1489 a_6122_3184.t4 a_6027_3169.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1454 a_6122_1457.t1 a_6027_1442.t3 VDD.t1626 VDD.t1625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1455 a_4745_n4470.t1 SAEN.t24 a_4942_n4114.t0 VSS.t296 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1456 a_3833_n953.t10 WWL[12].t10 a_3822_693.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1457 a_7283_n953.t3 WWLD[5].t15 a_7272_n512.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1458 VDD.t802 a_8422_4686.t3 a_8327_4671.t1 VDD.t801 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1459 a_7752_960.t0 WWL[11].t11 a_8020_4887.t26 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1460 a_402_n1770.t1 SA_OUT[0].t3 a_310_n1371.t1 VSS.t1902 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1461 a_8433_n953.t9 WWL[10].t7 a_8422_1216.t1 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1462 a_9218_n2086.t0 a_8977_n2234.t3 VSS.t2361 VSS.t2360 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1463 a_8792_4148.t0 VSS.t683 a_8340_n953.t13 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1464 a_6122_211.t0 a_6027_196.t3 VSS.t1151 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1465 a_372_2943.t2 a_277_2928.t3 VDD.t446 VDD.t445 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1466 VSS.t2159 a_2672_2943.t4 a_3042_2943.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1467 a_2577_4133.t0 WWLD[2].t8 a_2845_4887.t11 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1468 a_383_n953.t26 WWL[0].t7 a_372_3666.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1469 a_1892_2943.t0 RWLB[3].t1 a_1440_n953.t34 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1470 a_958_n953.t4 WWL[10].t8 a_947_1216.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1471 VSS.t2281 a_4397_693.t3 a_4767_693.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1472 a_8915_n30.t0 a_8902_n45.t3 VSS.t2476 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1473 a_7109_n4470.t0 SAEN.t25 a_7306_n4114.t0 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1474 a_1522_4445.t2 a_1427_4430.t3 VDD.t751 VDD.t750 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1475 a_3822_3907.t1 a_3727_3892.t4 VSS.t2440 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1476 VSS.t1071 a_4397_2421.t5 a_4302_2406.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1477 a_4315_1216.t0 a_4302_1201.t4 VSS.t105 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1478 a_3810_n1770.t1 PRE_VLSA.t15 VSS.t122 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1479 a_2097_n30.t1 a_2002_n45.t3 VDD.t1000 VDD.t999 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1480 VSS.t1260 a_6122_211.t3 a_6492_211.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1481 a_5547_1216.t1 a_5452_1201.t3 VDD.t761 VDD.t760 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1482 a_865_n1053.t1 a_852_n1068.t4 VSS.t1966 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1483 a_5452_n827.t0 WWLD[6].t13 a_5720_4887.t15 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1484 a_7642_452.t0 RWLB[13].t4 a_7190_n953.t22 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1485 a_372_n512.t1 a_277_n527.t4 VSS.t2265 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1486 a_13864_n8583.t1 ADC15_OUT[3].t3 a_13934_n8071.t2 VSS.t1443 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1487 a_742_n812.t0 VSS.t682 a_290_n953.t13 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1488 a_2108_n953.t1 WWL[2].t7 a_2097_3184.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1489 a_5547_1698.t1 a_5452_1683.t4 VSS.t1482 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1490 VSS.t2157 a_6697_4148.t4 a_6602_4133.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1491 a_8997_3907.t1 a_8902_3892.t5 VDD.t928 VDD.t927 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1492 a_8340_n953.t28 RWL[7].t4 a_8340_1939.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1493 a_865_n953.t27 RWL[7].t5 a_865_1939.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1494 a_2097_1216.t1 a_2002_1201.t5 VSS.t447 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1495 a_4883_n8071.t0 VCLP.t31 a_4745_n8071.t1 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1496 a_1317_1939.t1 RWLB[7].t3 a_865_n953.t31 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1497 a_8792_n1053.t0 VSS.t681 a_8340_n953.t7 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1498 VSS.t1857 a_4397_1939.t3 a_4767_1939.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1499 a_n3792_n6503.t1 VCLP.t32 a_n3827_n6849.t0 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1500 a_11776_n5850.t2 ADC13_OUT[1].t3 VDD.t509 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1501 a_4877_2647.t2 WWL[4].t7 a_5145_4887.t8 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1502 a_2015_n953.t39 RWL[13].t3 a_2015_452.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1503 a_n1233_n8583.t0 PRE_CLSA.t40 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1504 a_4448_n3770.t1 VCLP.t33 a_4413_n4116.t0 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1505 a_8340_1698.t1 a_8327_1683.t4 VSS.t1039 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 VSS.t85 a_947_452.t4 a_852_437.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1507 a_9008_n953.t20 WWLD[0].t10 a_8997_4686.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1508 VSS.t1793 a_4972_1939.t4 a_4877_1924.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1509 a_7247_n8071.t0 VCLP.t34 a_7109_n8071.t1 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1510 VDD.t664 a_1129_n8583.t3 ADC4_OUT[3].t1 VDD.t663 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1511 VDD.t1200 PRE_A.t3 a_8568_n2426.t3 VDD.t1199 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1512 a_1533_n953.t0 WWL[3].t6 a_1522_2943.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1513 VDD.t1499 a_947_2662.t4 a_852_2647.t0 VDD.t1498 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1514 a_865_1698.t0 a_852_1683.t5 VSS.t1591 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1515 a_4302_n527.t2 WWLD[5].t16 a_4570_4887.t5 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1516 a_3822_3425.t1 a_3727_3410.t4 VSS.t2497 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1517 a_4972_1457.t2 a_4877_1442.t3 VSS.t2211 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1518 VDD.t1591 a_n1233_n5850.t3 ADC2_OUT[1].t1 VDD.t1590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1519 a_3740_n953.t39 RWL[13].t4 a_3740_452.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1520 a_3617_3666.t0 RWLB[0].t4 a_3165_n953.t27 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1521 VSS.t2062 a_4972_2662.t4 a_5342_2662.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1522 a_4767_1698.t0 RWLB[8].t8 a_4315_n953.t27 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1523 a_3740_4686.t1 a_3727_4671.t4 VSS.t1602 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1524 VSS.t848 a_2672_452.t3 a_2577_437.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1525 a_6122_4686.t1 a_6027_4671.t3 VDD.t668 VDD.t667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1526 VSS.t1976 a_8997_2662.t5 a_8902_2647.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1527 VSS.t1577 a_867_n4378.t5 a_867_n4116.t1 VSS.t1573 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1528 a_7067_n30.t1 RWLB[15].t4 a_6615_n953.t39 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1529 a_8433_n953.t24 WWLD[1].t7 a_8422_4445.t1 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1530 a_8997_3425.t2 a_8902_3410.t5 VDD.t1065 VDD.t1064 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1531 a_5547_1216.t2 a_5452_1201.t4 VSS.t1563 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1532 VDD.t517 a_3822_2421.t4 a_3727_2406.t1 VDD.t516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1533 VDD.t1697 a_6122_2943.t3 a_6027_2928.t1 VDD.t1696 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1534 a_8327_2647.t1 WWL[4].t8 a_8595_4887.t10 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1535 a_958_n953.t18 WWLD[1].t8 a_947_4445.t1 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1536 a_8902_2165.t0 WWL[6].t9 a_9170_4887.t15 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1537 a_8792_n30.t0 RWLB[15].t5 a_8340_n953.t33 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1538 a_4315_4445.t1 a_4302_4430.t4 VSS.t2422 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1539 a_7752_4133.t2 WWLD[2].t9 a_8020_4887.t10 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1540 a_7067_2943.t1 RWLB[3].t2 a_6615_n953.t38 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1541 a_3152_960.t0 WWL[11].t12 a_3420_4887.t4 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1542 a_8902_437.t2 WWL[13].t7 a_9170_4887.t21 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1543 a_1522_211.t0 a_1427_196.t3 VSS.t1894 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1544 a_852_2928.t0 WWL[3].t7 a_1120_4887.t14 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1545 a_4890_n953.t11 VSS.t680 a_4890_3907.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1546 VSS.t823 a_8422_2421.t4 a_8327_2406.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1547 VDD.t1716 a_4972_2180.t3 a_4877_2165.t1 VDD.t1715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1548 a_6122_1939.t1 a_6027_1924.t4 VSS.t976 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1549 a_5547_4445.t0 a_5452_4430.t3 VDD.t542 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1550 a_8340_1216.t0 a_8327_1201.t4 VSS.t504 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1551 a_1317_452.t0 RWLB[13].t5 a_865_n953.t23 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1552 a_2590_n953.t24 RWL[11].t2 a_2590_975.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1553 a_6697_975.t1 a_6602_960.t4 VSS.t94 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1554 a_290_3666.t1 a_277_3651.t4 VSS.t2203 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1555 VSS.t2072 a_8997_2180.t3 a_9367_2180.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1556 a_865_1216.t0 a_852_1201.t5 VSS.t1478 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1557 a_7260_n1770.t0 a_7445_4887.t27 a_7453_n1770.t1 VSS.t2400 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1558 VSS.t1265 a_7847_4148.t3 a_8217_4148.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1559 VSS.t1286 a_1522_211.t3 a_1892_211.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1560 SA_OUT[1].t0 PRE_VLSA.t16 VDD.t1145 VDD.t1144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1561 a_4192_3666.t1 RWLB[0].t5 a_3740_n953.t28 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1562 a_4767_1216.t1 RWLB[10].t8 a_4315_n953.t35 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1563 a_3833_n953.t24 WWL[4].t9 a_3822_2662.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1564 a_1440_n953.t8 VSS.t679 a_1440_n512.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1565 a_7039_n7216.t1 ADC9_OUT[2].t3 VDD.t1712 VDD.t1673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1566 a_n3357_n8071.t1 Iref3.t5 a_n3298_n8026.t1 VSS.t824 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1567 a_3258_n953.t11 WWLD[2].t10 a_3247_4148.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1568 a_6133_n953.t24 WWL[2].t8 a_6122_3184.t1 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1569 a_2097_4445.t0 a_2002_4430.t5 VSS.t1093 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1570 VSS.t1990 a_1522_3907.t4 a_1427_3892.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1571 a_5465_n953.t28 RWL[0].t9 a_5465_3666.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1572 a_8422_3666.t0 a_8327_3651.t4 VSS.t1271 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1573 a_7190_975.t1 a_7177_960.t4 VSS.t2035 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1574 a_8217_3907.t0 VSS.t678 a_7765_n953.t11 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1575 VDD.t1612 a_4397_1939.t4 a_4302_1924.t2 VDD.t1611 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1576 a_947_3666.t1 a_852_3651.t4 VSS.t1391 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1577 a_2015_3184.t1 a_2002_3169.t4 VSS.t2325 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1578 a_5342_1939.t1 RWLB[7].t4 a_4890_n953.t40 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1579 VSS.t1969 a_8422_1939.t4 a_8792_1939.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1580 a_3247_3184.t0 a_3152_3169.t3 VDD.t355 VDD.t354 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1581 a_4408_n953.t3 WWL[5].t6 a_4397_2421.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1582 a_8422_n30.t1 a_8327_n45.t4 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1583 a_4890_n953.t5 VSS.t677 a_4890_n271.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1584 SA_OUT[6].t2 PRE_VLSA.t17 VDD.t1143 VDD.t1142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1585 a_277_n1068.t2 WWLD[7].t9 a_545_4887.t26 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1586 a_4972_4686.t1 a_4877_4671.t3 VSS.t2286 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1587 a_902_n8026.t1 VCLP.t35 a_867_n7825.t0 VSS.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1588 VSS.t1991 a_2097_3666.t5 a_2002_3651.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1589 VDD.t906 a_8422_2662.t3 a_8327_2647.t0 VDD.t905 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1590 VSS.t299 SAEN.t26 a_9178_n8026.t0 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1591 a_8221_n4483.t2 ADC10_OUT[0].t4 VDD.t1511 VDD.t1510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1592 a_4890_n953.t21 RWL[1].t3 a_4890_3425.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1593 a_8792_1698.t0 RWLB[8].t9 a_8340_n953.t29 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1594 a_7642_3666.t1 RWLB[0].t6 a_7190_n953.t25 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1595 VSS.t1496 a_5632_n6430# a_11549_n6503.t0 VSS.t281 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1596 VSS.t300 SAEN.t27 a_n3792_n5293.t0 VSS.t277 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1597 a_1427_3651.t2 WWL[0].t8 a_1695_4887.t26 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1598 a_1522_2421.t2 a_1427_2406.t3 VDD.t1849 VDD.t1848 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1599 a_2577_1683.t2 WWL[8].t8 a_2845_4887.t10 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1600 VSS.t1779 a_1522_n271.t4 a_1427_n286.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1601 a_11776_n5850.t0 PRE_CLSA.t41 VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1602 VSS.t2169 a_3247_n1053.t3 a_3617_n1053.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1603 a_5547_4445.t1 a_5452_4430.t4 VSS.t898 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1604 a_6708_n953.t16 WWLD[2].t11 a_6697_4148.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1605 a_7858_n953.t20 WWL[6].t10 a_7847_2180.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1606 a_8422_975.t0 a_8327_960.t3 VSS.t2183 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1607 a_1522_n271.t1 a_1427_n286.t3 VDD.t1847 VDD.t1846 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1608 a_8410_n1770.t2 a_8595_4887.t27 a_8603_n1770.t1 VSS.t2192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1609 a_8915_n953.t29 RWL[0].t10 a_8915_3666.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1610 SA_OUT[3].t0 PRE_VLSA.t18 VDD.t1141 VDD.t1140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1611 VSS.t1882 a_2672_975.t3 a_2577_960.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1612 a_2467_n30.t0 RWLB[15].t6 a_2015_n953.t34 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1613 VSS.t2067 a_6677_n2234.t3 a_6800_n2132.t0 VSS.t2066 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1614 VSS.t1914 a_1522_3425.t4 a_1427_3410.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1615 a_383_n953.t22 WWL[15].t10 a_372_n30.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1616 a_9367_1457.t1 RWLB[9].t3 a_8915_n953.t39 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1617 a_n1163_n8071.t0 SAEN.t28 a_n966_n8026.t0 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1618 a_14072_n5338.t0 VCLP.t36 a_13934_n5338.t1 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1619 a_n3792_n3770.t1 VCLP.t37 a_n3827_n4116.t0 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1620 a_8217_3425.t1 RWLB[1].t1 a_7765_n953.t34 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1621 a_3822_4148.t0 a_3727_4133.t3 VDD.t690 VDD.t689 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1622 a_6697_3184.t2 a_6602_3169.t3 VDD.t918 VDD.t917 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1623 a_3152_1442.t0 WWL[9].t11 a_3420_4887.t21 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1624 VDD.t171 PRE_CLSA.t42 ADC13_OUT[0].t0 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1625 a_8340_4445.t1 a_8327_4430.t4 VSS.t1572 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1626 VSS.t1076 a_6697_1698.t4 a_6602_1683.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1627 VSS.t303 SAEN.t29 a_n2642_n8026.t0 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1628 VSS.t1657 a_5547_3666.t5 a_5452_3651.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1629 a_4877_2928.t0 WWL[3].t8 a_5145_4887.t7 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1630 a_4302_437.t1 WWL[13].t8 a_4570_4887.t19 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1631 a_865_4445.t1 a_852_4430.t5 VSS.t2415 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1632 VDD.t1823 a_8997_2180.t4 a_8902_2165.t1 VDD.t1822 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1633 a_277_196.t0 WWL[14].t13 a_545_4887.t11 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1634 VDD.t898 a_7847_4148.t4 a_7752_4133.t0 VDD.t897 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1635 a_6040_n953.t0 RWL[15].t3 a_6040_n30.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1636 SA_OUT[8].t0 PRE_VLSA.t19 VDD.t1139 VDD.t1138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1637 a_947_n1053.t1 a_852_n1068.t5 VDD.t1726 VDD.t1725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1638 VSS.t1618 a_6697_n812.t4 a_6602_n827.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1639 a_4767_4445.t1 VSS.t676 a_4315_n953.t18 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1640 VDD.t1577 a_372_4148.t3 a_277_4133.t2 VDD.t1576 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1641 VSS.t1024 a_n2677_n4378.t6 a_n2677_n7825.t1 VSS.t1021 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1642 VSS.t1891 a_2672_3907.t4 a_3042_3907.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1643 VSS.t2073 a_3247_1457.t3 a_3617_1457.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1644 a_3247_3184.t2 a_3152_3169.t4 VSS.t1275 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1645 a_9008_n953.t12 WWL[4].t10 a_8997_2662.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1646 a_290_n953.t16 VSS.t675 a_290_n1053.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1647 a_8792_1216.t1 RWLB[10].t9 a_8340_n953.t34 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1648 a_2577_1201.t0 WWL[10].t9 a_2845_4887.t2 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1649 a_5558_n953.t15 WWL[14].t14 a_5547_211.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1650 VSS.t2425 a_3822_n1053.t3 a_4192_n1053.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1651 a_7283_n953.t16 WWLD[2].t12 a_7272_4148.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1652 a_11984_n8071.t1 Iref3.t6 a_12043_n8026.t1 VSS.t825 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1653 VDD.t1091 a_1522_3666.t3 a_1427_3651.t0 VDD.t1090 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1654 a_3740_2662.t0 a_3727_2647.t4 VSS.t775 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1655 a_2590_975.t1 a_2577_960.t4 VSS.t1737 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1656 a_3165_4148.t1 a_3152_4133.t5 VSS.t854 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1657 a_6027_3892.t2 WWLD[3].t9 a_6295_4887.t8 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1658 a_6040_3184.t0 a_6027_3169.t4 VSS.t432 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1659 a_6122_2662.t1 a_6027_2647.t3 VDD.t1310 VDD.t1309 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1660 a_7847_211.t0 a_7752_196.t3 VSS.t1331 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1661 VSS.t1772 a_1522_n512.t4 a_1892_n512.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1662 a_5857_n5850.t2 ADC8_OUT[1].t3 VDD.t1089 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1663 a_6602_1924.t0 WWL[7].t11 a_6870_4887.t16 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1664 a_8327_2928.t0 WWL[3].t9 a_8595_4887.t9 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 a_8433_n953.t6 WWL[5].t7 a_8422_2421.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1666 VDD.t173 PRE_CLSA.t43 ADC4_OUT[1].t0 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1667 a_6615_693.t0 a_6602_678.t4 VSS.t1099 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 a_2097_n512.t1 a_2002_n527.t3 VDD.t1756 VDD.t1755 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1669 VSS.t2114 a_6122_3666.t4 a_6027_3651.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1670 a_2467_3184.t1 RWLB[2].t7 a_2015_n953.t44 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1671 VSS.t1029 a_6697_1216.t4 a_6602_1201.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1672 VDD.t1956 a_3822_n30.t3 a_3727_n45.t2 VDD.t1955 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1673 a_3822_n30.t2 a_3727_n45.t4 VDD.t1962 VDD.t1961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1674 a_1337_n8071.t1 Iref3.t7 a_1396_n8026.t1 VSS.t826 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1675 a_2311_n8583.t0 PRE_CLSA.t44 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1676 a_958_n953.t2 WWL[5].t8 a_947_2421.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1677 VSS.t1183 a_2672_n271.t4 a_3042_n271.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1678 a_5053_n2086.t1 WE.t13 a_4983_n953.t13 VSS.t2386 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1679 a_4315_2421.t0 a_4302_2406.t4 VSS.t1094 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1680 a_1522_2180.t1 a_1427_2165.t4 VSS.t1639 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1681 a_290_n953.t19 RWL[9].t2 a_290_1457.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1682 VDD.t1922 a_3247_n1053.t4 a_3152_n1068.t0 VDD.t1921 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1683 a_7752_1683.t2 WWL[8].t9 a_8020_4887.t11 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1684 a_6027_437.t2 WWL[13].t9 a_6295_4887.t17 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1685 a_7283_n953.t23 WWL[13].t10 a_7272_452.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1686 a_8340_211.t1 a_8327_196.t4 VSS.t1907 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1687 a_4315_n271.t1 a_4302_n286.t4 VSS.t1084 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1688 a_9405_n8583.t1 ADC11_OUT[3].t3 VDD.t1851 VDD.t1850 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1689 a_4890_n812.t1 a_4877_n827.t5 VSS.t226 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1690 a_2097_n1053.t2 a_2002_n1068.t4 VDD.t540 VDD.t539 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1691 a_1522_n1053.t0 a_1427_n1068.t4 VSS.t2452 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1692 a_7272_n812.t1 a_7177_n827.t3 VDD.t1475 VDD.t1474 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1693 VSS.t1554 a_2672_3425.t4 a_3042_3425.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1694 a_5547_2421.t0 a_5452_2406.t3 VDD.t759 VDD.t758 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1695 VSS.t875 a_3822_1457.t3 a_4192_1457.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1696 VSS.t1705 a_7272_n1053.t4 a_7642_n1053.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1697 a_1533_n953.t9 WWLD[3].t10 a_1522_3907.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1698 VSS.t2518 a_7847_975.t5 a_7752_960.t2 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1699 a_1440_n953.t37 EN.t3 a_n1495_n4378.t3 VSS.t2044 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1700 a_3822_975.t0 a_3727_960.t3 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1701 VDD.t1364 a_4972_693.t4 a_4877_678.t1 VDD.t1363 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1702 a_5547_n271.t0 a_5452_n286.t3 VDD.t771 VDD.t770 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1703 a_9367_4686.t0 VSS.t674 a_8915_n953.t15 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1704 a_7765_2180.t1 a_7752_2165.t5 VSS.t1671 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1705 VSS.t1141 a_7847_1698.t3 a_8217_1698.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1706 a_7190_n953.t42 RWL[12].t5 a_7190_693.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1707 a_2683_n953.t26 WWLD[7].t10 a_2672_n1053.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1708 a_3152_4671.t2 WWLD[0].t11 a_3420_4887.t7 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1709 a_6615_4148.t1 a_6602_4133.t4 VSS.t1096 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1710 VSS.t1194 a_372_n1053.t4 a_277_n1068.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1711 a_2097_2421.t0 a_2002_2406.t5 VSS.t1781 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1712 VSS.t1014 a_6122_693.t4 a_6027_678.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1713 VDD.t702 a_6697_693.t4 a_6602_678.t1 VDD.t701 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1714 a_7847_4148.t2 a_7752_4133.t3 VDD.t978 VDD.t977 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1715 a_6027_3410.t0 WWL[1].t10 a_6295_4887.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1716 a_3258_n953.t12 WWL[8].t10 a_3247_1698.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1717 a_7177_1442.t2 WWL[9].t12 a_7445_4887.t15 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1718 VSS.t2085 a_7847_n812.t3 a_8217_n812.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1719 a_2108_n953.t26 WWL[0].t9 a_2097_3666.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1720 a_2097_n271.t0 a_2002_n286.t5 VSS.t2150 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1721 a_5917_3184.t0 RWLB[2].t8 a_5465_n953.t46 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1722 VSS.t1333 a_7847_211.t3 a_8217_211.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1723 VSS.t794 a_3247_4686.t3 a_3617_4686.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1724 VDD.t456 a_6122_3907.t3 a_6027_3892.t0 VDD.t455 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1725 VDD.t1821 a_3247_1457.t4 a_3152_1442.t1 VDD.t1820 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1726 a_1168_n2086.t0 a_927_n2234.t3 VSS.t2513 VSS.t2512 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1727 a_3258_n953.t7 WWLD[6].t14 a_3247_n812.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1728 a_3266_n8026.t1 VCLP.t38 a_3231_n7825.t0 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1729 VDD.t1291 a_12963_n8583.t3 ADC14_OUT[3].t1 VDD.t1290 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1730 VSS.t986 a_6693_n2422.t5 a_9143_n4116.t1 VSS.t982 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1731 a_8792_4445.t1 VSS.t673 a_8340_n953.t17 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1732 VSS.t305 SAEN.t30 a_11549_n3770.t0 VSS.t304 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1733 a_4972_2662.t1 a_4877_2647.t3 VSS.t838 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1734 VSS.t1612 a_7272_1457.t4 a_7642_1457.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1735 a_1533_n953.t16 WWLD[4].t8 a_1522_n271.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1736 VDD.t1019 a_9405_n4483.t4 ADC11_OUT[0].t2 VDD.t1018 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1737 a_2577_4430.t2 WWLD[1].t9 a_2845_4887.t15 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1738 a_4397_4148.t1 a_4302_4133.t5 VSS.t1818 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1739 a_7272_3184.t1 a_7177_3169.t4 VSS.t1465 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1740 a_7752_1201.t2 WWL[10].t10 a_8020_4887.t4 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1741 VSS.t1732 a_2775_n2132.t2 a_2753_n2086.t1 VSS.t1731 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 VSS.t1065 a_3231_n4378.t4 a_3231_n6849.t1 VSS.t1064 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1743 a_1533_n953.t2 WWL[1].t11 a_1522_3425.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1744 a_2683_n953.t12 WWL[9].t13 a_2672_1457.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 VSS.t1697 a_372_1457.t4 a_277_1442.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1746 a_2590_n953.t35 EN.t4 a_867_n4378.t2 VSS.t1944 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1747 VSS.t2254 a_6697_n512.t5 a_7067_n512.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1748 a_7190_4148.t1 a_7177_4133.t4 VSS.t1059 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1749 a_5547_2421.t1 a_5452_2406.t4 VSS.t1132 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1750 VSS.t792 a_7847_1216.t3 a_8217_1216.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1751 VSS.t1057 a_372_452.t4 a_277_437.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1752 a_7177_n45.t0 WWL[15].t11 a_7445_4887.t11 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1753 a_6708_n953.t15 WWL[8].t11 a_6697_1698.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1754 a_5547_n271.t1 a_5452_n286.t4 VSS.t1143 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1755 VSS.t1711 a_6697_4445.t4 a_6602_4430.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1756 a_6492_693.t0 RWLB[12].t2 a_6040_n953.t19 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1757 VDD.t648 a_6122_n271.t3 a_6027_n286.t0 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1758 VSS.t1925 a_n314_n4378.t4 a_n314_n6849.t1 VSS.t1924 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1759 a_2084_n6503.t2 a_2311_n7216.t4 ADC5_OUT[2].t1 VSS.t1106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1760 a_3258_n953.t3 WWL[10].t11 a_3247_1216.t1 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1761 a_2015_211.t1 a_2002_196.t4 VSS.t1257 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1762 a_290_n953.t3 VSS.t672 a_290_4686.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1763 VDD.t1636 a_7272_975.t3 a_7177_960.t2 VDD.t1635 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1764 a_6708_n953.t10 WWLD[6].t15 a_6697_n812.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1765 a_6492_3184.t1 RWLB[2].t9 a_6040_n953.t31 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1766 a_1317_n512.t0 VSS.t671 a_865_n953.t5 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1767 VDD.t1137 PRE_VLSA.t20 a_3760_n1371.t2 VDD.t1136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1768 VSS.t1388 a_3822_4686.t3 a_4192_4686.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1769 VDD.t773 a_6122_3425.t3 a_6027_3410.t1 VDD.t772 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1770 a_8340_2421.t1 a_8327_2406.t4 VSS.t2004 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1771 a_8997_2180.t0 a_8902_2165.t4 VSS.t1860 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1772 VSS.t1495 a_5632_n6430# a_5630_n6503.t0 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1773 a_8402_n2234.t0 Din[14].t1 VSS.t1714 VSS.t1713 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1774 a_1440_n953.t6 VSS.t670 a_1440_4148.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1775 a_7847_4148.t1 a_7752_4133.t4 VSS.t1338 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1776 a_7765_n953.t30 RWL[2].t10 a_7765_3184.t1 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1777 a_2590_n953.t32 RWL[6].t3 a_2590_2180.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1778 a_3822_1698.t1 a_3727_1683.t3 VDD.t1896 VDD.t1895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1779 a_3247_452.t1 a_3152_437.t3 VSS.t2052 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1780 a_1427_437.t2 WWL[13].t11 a_1695_4887.t20 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 a_3740_211.t1 a_3727_196.t4 VSS.t1186 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1782 a_8340_n271.t1 a_8327_n286.t4 VSS.t1297 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1783 a_5857_n5850.t0 PRE_CLSA.t45 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1784 a_2318_n2086.t1 a_2077_n2234.t3 VSS.t1784 VSS.t1783 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1785 a_865_2421.t1 a_852_2406.t5 VSS.t2283 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1786 a_2683_n953.t24 WWL[13].t12 a_2672_452.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1787 a_6295_4887.t4 PRE_SRAM.t16 VDD.t2041 VDD.t2040 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1788 VSS.t1588 a_372_975.t4 a_742_975.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1789 a_865_n271.t1 a_852_n286.t5 VSS.t1570 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1790 a_3042_n812.t0 VSS.t669 a_2590_n953.t5 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1791 a_4767_2421.t0 RWLB[5].t9 a_4315_n953.t40 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1792 VDD.t769 a_7847_1698.t4 a_7752_1683.t0 VDD.t768 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1793 a_n2207_n7203.t0 VCLP.t39 a_n2345_n7203.t1 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1794 VSS.t1494 a_5632_n6430# a_7994_n6503.t0 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1795 VSS.t950 a_3925_n2132.t2 a_3903_n2086.t1 VSS.t949 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1796 VDD.t1240 a_372_1698.t3 a_277_1683.t1 VDD.t1239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1797 a_4972_452.t0 a_4877_437.t3 VSS.t1545 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1798 a_4767_n271.t0 VSS.t668 a_4315_n953.t6 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1799 a_7177_4671.t0 WWLD[0].t12 a_7445_4887.t20 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1800 a_1440_3907.t1 a_1427_3892.t4 VSS.t2110 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1801 a_2590_n953.t42 RWL[12].t6 a_2590_693.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1802 VDD.t179 PRE_CLSA.t46 ADC11_OUT[0].t0 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1803 VDD.t1841 a_7847_n812.t4 a_7752_n827.t2 VDD.t1840 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1804 VSS.t1906 a_4397_3184.t5 a_4302_3169.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1805 a_3165_n953.t30 RWL[7].t6 a_3165_1939.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1806 VDD.t1780 a_2097_211.t4 a_2002_196.t2 VDD.t1779 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1807 VDD.t181 PRE_CLSA.t47 ADC8_OUT[0].t0 VDD.t180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1808 VDD.t1135 PRE_VLSA.t21 a_6635_n1371.t0 VDD.t1134 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1809 a_3740_2943.t1 a_3727_2928.t4 VSS.t1631 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1810 a_742_452.t1 RWLB[13].t6 a_290_n953.t21 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1811 a_5558_n953.t11 WWLD[5].t17 a_5547_n512.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1812 a_6122_2943.t2 a_6027_2928.t3 VDD.t484 VDD.t483 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1813 a_947_1939.t0 a_852_1924.t3 VDD.t379 VDD.t378 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1814 VSS.t1295 a_1522_693.t4 a_1427_678.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1815 VDD.t558 a_372_n812.t3 a_277_n827.t1 VDD.t557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 VDD.t464 a_3247_4686.t4 a_3152_4671.t0 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1817 a_6133_n953.t25 WWL[0].t10 a_6122_3666.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1818 a_7283_n953.t17 WWL[8].t12 a_7272_1698.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1819 a_6708_n953.t3 WWL[10].t12 a_6697_1216.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1820 a_6122_693.t2 a_6027_678.t4 VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 VDD.t1202 PRE_A.t4 a_2049_n4378.t2 VDD.t1201 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1822 VSS.t481 a_947_2943.t3 a_1317_2943.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1823 VSS.t919 a_7272_4686.t4 a_7642_4686.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1824 VSS.t1599 a_3247_211.t3 a_3617_211.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1825 a_10589_n5850.t2 ADC12_OUT[1].t3 VDD.t1296 VDD.t1276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1826 a_935_n1770.t1 PRE_VLSA.t22 VSS.t118 VSS.t117 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1827 a_2015_3666.t1 a_2002_3651.t4 VSS.t1794 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 a_3165_1698.t1 a_3152_1683.t5 VSS.t1652 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1829 a_3701_n8071.t1 Iref3.t8 a_3760_n8026.t1 VSS.t827 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1830 a_7283_n953.t11 WWLD[6].t16 a_7272_n812.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1831 a_7752_4430.t2 WWLD[1].t10 a_8020_4887.t15 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1832 a_1892_n1053.t1 VSS.t667 a_1440_n953.t3 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1833 a_7847_693.t1 a_7752_678.t4 VDD.t968 VDD.t967 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1834 VDD.t1133 PRE_VLSA.t23 a_4910_n1371.t2 VDD.t1132 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1835 a_2683_n953.t20 WWLD[0].t13 a_2672_4686.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1836 a_3247_3666.t0 a_3152_3651.t3 VDD.t2148 VDD.t2147 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1837 a_3822_1216.t1 a_3727_1201.t3 VDD.t1473 VDD.t1472 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1838 VDD.t183 PRE_CLSA.t48 ADC1_OUT[0].t0 VDD.t182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1839 a_6122_n512.t1 a_6027_n527.t4 VSS.t1457 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1840 VSS.t1292 a_372_4686.t4 a_277_4671.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1841 a_6065_n8071.t1 Iref3.t9 a_6124_n8026.t1 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1842 a_852_n45.t0 WWL[15].t12 a_1120_4887.t18 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1843 VDD.t1204 PRE_A.t5 a_n1495_n4378.t2 VDD.t1203 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1844 VSS.t1307 a_7847_4445.t3 a_8217_4445.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1845 VDD.t462 a_7847_1216.t4 a_7752_1201.t0 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1846 VSS.t2081 a_2672_2180.t3 a_2577_2165.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1847 a_6615_n953.t32 RWL[7].t7 a_6615_1939.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1848 VSS.t1212 a_5543_n2422.t6 a_6777_n7825.t1 VSS.t1209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1849 a_2590_1457.t0 a_2577_1442.t4 VSS.t1299 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1850 VDD.t325 a_372_1216.t3 a_277_1201.t1 VDD.t324 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1851 a_4397_n30.t1 a_4302_n45.t4 VSS.t962 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1852 a_3258_n953.t16 WWLD[1].t11 a_3247_4445.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1853 a_1440_3425.t1 a_1427_3410.t4 VSS.t2038 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1854 a_4397_1939.t2 a_4302_1924.t3 VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1855 a_4972_1457.t1 a_4877_1442.t4 VDD.t1954 VDD.t1953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1856 a_2577_n45.t2 WWL[15].t13 a_2845_4887.t9 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1857 a_9367_2662.t1 RWLB[4].t3 a_8915_n953.t47 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1858 VSS.t1543 a_4972_452.t3 a_5342_452.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1859 a_372_n812.t1 a_277_n827.t4 VSS.t1078 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1860 a_1892_693.t0 RWLB[12].t3 a_1440_n953.t20 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1861 a_6152_n1770.t1 a_6133_n953.t27 a_6110_n1770.t2 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1862 VDD.t1131 PRE_VLSA.t24 a_7785_n1371.t0 VDD.t1130 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1863 a_2845_4887.t19 PRE_SRAM.t17 a_2683_n953.t21 VDD.t2042 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1864 a_3152_2647.t2 WWL[4].t11 a_3420_4887.t24 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1865 a_7283_n953.t4 WWL[10].t13 a_7272_1216.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1866 a_6615_1698.t1 a_6602_1683.t4 VSS.t1935 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1867 VSS.t1317 a_3247_1939.t5 a_3152_1924.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1868 a_5342_n512.t0 VSS.t666 a_4890_n953.t8 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1869 a_1337_n5338.t0 VCLP.t40 a_1199_n5338.t1 VSS.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1870 VDD.t1206 PRE_A.t6 a_4393_n2422.t2 VDD.t1205 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1871 a_2672_3907.t1 a_2577_3892.t4 VSS.t1892 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1872 a_7847_1698.t2 a_7752_1683.t3 VDD.t1853 VDD.t1852 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1873 a_3165_1216.t0 a_3152_1201.t5 VSS.t998 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1874 a_865_n953.t33 EN.t5 a_n2677_n4378.t2 VSS.t1945 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1875 a_6697_3666.t1 a_6602_3651.t3 VDD.t1258 VDD.t1257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1876 VSS.t92 a_n3827_n4378.t5 a_n3827_n5092.t1 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1877 VDD.t1768 a_3822_3184.t4 a_3727_3169.t2 VDD.t1767 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1878 a_4972_2943.t1 a_4877_2928.t3 VSS.t929 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1879 VSS.t1372 a_3247_2662.t3 a_3617_2662.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1880 VSS.t101 a_4393_n2422.t5 a_4413_n5092.t1 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1881 a_7847_n1053.t0 a_7752_n1068.t4 VDD.t785 VDD.t784 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1882 a_11776_n5850.t1 ADC13_OUT[1].t4 a_11846_n5338.t2 VSS.t862 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1883 a_8792_2421.t1 RWLB[5].t10 a_8340_n953.t42 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1884 a_4302_n827.t2 WWLD[6].t17 a_4570_4887.t7 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1885 VSS.t1413 a_1522_4148.t4 a_1892_4148.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1886 a_2577_2406.t2 WWL[5].t9 a_2845_4887.t4 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1887 a_8792_n271.t0 VSS.t665 a_8340_n953.t12 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1888 a_3493_n7216.t1 ADC6_OUT[2].t3 VDD.t1055 VDD.t1054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1889 VDD.t185 PRE_CLSA.t49 ADC0_OUT[0].t0 VDD.t184 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1890 a_9027_n1770.t1 a_9008_n953.t27 a_8985_n1770.t1 VSS.t2164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1891 a_4397_1698.t1 a_4302_1683.t5 VSS.t2342 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1892 a_5917_n30.t1 RWLB[15].t7 a_5465_n953.t37 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1893 a_2577_n286.t0 WWLD[4].t9 a_2845_4887.t16 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1894 a_6708_n953.t17 WWLD[1].t12 a_6697_4445.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1895 a_3247_3666.t1 a_3152_3651.t4 VSS.t2340 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1896 VSS.t242 a_8422_3184.t4 a_8327_3169.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1897 a_7190_n953.t26 RWL[7].t8 a_7190_1939.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1898 a_8422_1457.t1 a_8327_1442.t3 VDD.t732 VDD.t731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1899 VDD.t1208 PRE_A.t7 a_867_n4378.t3 VDD.t1207 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1900 a_n1460_n5293.t2 a_n1233_n5850.t4 ADC2_OUT[1].t2 VSS.t1837 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1901 a_2084_n3770.t2 a_2311_n4483.t3 ADC5_OUT[0].t2 VSS.t458 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1902 VDD.t416 a_947_2943.t4 a_852_2928.t1 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1903 a_372_3907.t1 a_277_3892.t3 VDD.t1992 VDD.t1991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1904 a_1892_3907.t0 VSS.t664 a_1440_n953.t13 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1905 a_3727_2165.t2 WWL[6].t11 a_3995_4887.t11 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1906 a_290_975.t1 a_277_960.t4 VSS.t1221 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1907 a_1522_693.t2 a_1427_678.t4 VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1908 a_6122_n30.t1 a_6027_n45.t3 VSS.t1750 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1909 a_4448_n6503.t1 a_4675_n7216.t4 ADC7_OUT[2].t2 VSS.t1449 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1910 SA_OUT[4].t0 a_2610_n1371.t3 VDD.t742 VDD.t741 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1911 VSS.t927 a_4972_2943.t4 a_5342_2943.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1912 VSS.t307 SAEN.t31 a_5630_n3770.t0 VSS.t306 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1913 VSS.t502 a_6697_2421.t4 a_6602_2406.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1914 a_7190_1698.t1 a_7177_1683.t4 VSS.t2140 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1915 VSS.t1710 a_6122_n30.t5 a_6027_n45.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1916 a_3822_4445.t0 a_3727_4430.t3 VDD.t676 VDD.t675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1917 a_6040_3666.t1 a_6027_3651.t4 VSS.t1585 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1918 a_6615_1216.t1 a_6602_1201.t4 VSS.t1774 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1919 VDD.t187 PRE_CLSA.t50 ADC9_OUT[2].t0 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1920 a_13934_n8071.t0 SAEN.t32 a_14131_n8026.t0 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1921 VSS.t1411 a_8997_2943.t5 a_8902_2928.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1922 VSS.t1651 a_3822_1939.t4 a_3727_1924.t2 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1923 a_n2642_n8026.t1 VCLP.t41 a_n2677_n7825.t0 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1924 a_2015_n953.t15 VSS.t663 a_2015_n1053.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1925 a_290_n953.t46 RWL[4].t3 a_290_2662.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1926 a_3247_211.t1 a_3152_196.t4 VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1927 a_n1233_n5850.t0 PRE_CLSA.t51 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1928 a_4675_n4483.t1 ADC7_OUT[0].t4 VDD.t894 VDD.t893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1929 a_n52_n4483.t2 ADC3_OUT[0].t4 VDD.t1538 VDD.t1537 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1930 a_2672_3425.t1 a_2577_3410.t4 VSS.t241 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1931 a_7847_1216.t2 a_7752_1201.t3 VDD.t454 VDD.t453 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1932 a_3235_n1770.t0 a_3420_4887.t27 a_3428_n1770.t0 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1933 VDD.t944 a_7847_4445.t4 a_7752_4430.t0 VDD.t943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1934 a_13637_n8026.t1 VCLP.t42 a_13602_n7825.t0 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1935 VSS.t310 SAEN.t33 a_7994_n3770.t0 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1936 a_2467_3666.t0 RWLB[0].t7 a_2015_n953.t22 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1937 VSS.t1067 a_3822_2662.t3 a_4192_2662.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1938 a_4315_975.t1 a_4302_960.t4 VSS.t2107 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1939 VDD.t191 PRE_CLSA.t52 ADC3_OUT[3].t0 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1940 VDD.t1271 a_1129_n5850.t3 ADC4_OUT[1].t1 VDD.t1270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1941 a_n2207_n4470.t0 VCLP.t43 a_n2345_n4470.t1 VSS.t201 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1942 VSS.t1667 a_7847_2180.t5 a_7752_2165.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1943 VSS.t1493 a_5632_n6430# a_10362_n6503.t1 VSS.t289 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1944 a_2590_4686.t1 a_2577_4671.t4 VSS.t881 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1945 VDD.t1928 a_372_4445.t3 a_277_4430.t1 VDD.t1927 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1946 a_4408_n953.t26 WWL[2].t9 a_4397_3184.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1947 VDD.t896 a_8422_211.t4 a_8327_196.t2 VDD.t895 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 a_4972_4686.t2 a_4877_4671.t4 VDD.t2108 VDD.t2107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1949 a_1440_n953.t33 RWL[8].t6 a_1440_1698.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1950 a_7847_1698.t1 a_7752_1683.t4 VSS.t2092 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1951 VDD.t1059 a_2672_1939.t3 a_2577_1924.t1 VDD.t1058 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1952 VSS.t1397 a_8993_n2422.t4 a_13602_n6849.t1 VSS.t1396 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1953 a_8020_4887.t21 PRE_SRAM.t18 a_7858_n953.t25 VDD.t2043 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1954 a_4397_1216.t0 a_4302_1201.t5 VSS.t66 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1955 a_n3565_n7216.t2 ADC0_OUT[2].t4 a_n3495_n7203.t1 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1956 a_7283_n953.t18 WWLD[1].t13 a_7272_4445.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1957 a_1440_n953.t5 VSS.t662 a_1440_n812.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1958 a_3617_1939.t1 RWLB[7].t5 a_3165_n953.t25 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1959 a_1510_n1770.t2 a_1695_4887.t27 a_1703_n1770.t1 VSS.t1816 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1960 a_7177_2647.t2 WWL[4].t12 a_7445_4887.t10 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1961 a_6812_n8026.t2 a_7039_n8583.t4 ADC9_OUT[3].t1 VSS.t991 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1962 a_372_3425.t1 a_277_3410.t3 VDD.t1900 VDD.t1899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1963 a_1522_3184.t1 a_1427_3169.t3 VDD.t1746 VDD.t1745 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1964 VDD.t1308 a_n3565_n4483.t4 ADC0_OUT[0].t1 VDD.t1307 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1965 a_3165_4445.t1 a_3152_4430.t5 VSS.t2071 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1966 a_1892_3425.t1 RWLB[1].t2 a_1440_n953.t28 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1967 a_9008_n953.t24 WWL[13].t13 a_8997_452.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1968 VDD.t193 PRE_CLSA.t53 ADC12_OUT[0].t0 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1969 VSS.t2050 a_7272_1939.t4 a_7177_1924.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1970 a_2015_n953.t17 RWL[9].t3 a_2015_1457.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1971 a_6812_n6503.t2 a_5743_n6391# a_6777_n6849.t0 VSS.t178 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X1972 VDD.t1057 a_3247_2662.t4 a_3152_2647.t1 VDD.t1056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1973 a_6602_n527.t0 WWLD[5].t18 a_6870_4887.t12 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1974 a_3833_n953.t0 WWL[3].t10 a_3822_2943.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1975 a_7190_1216.t1 a_7177_1201.t4 VSS.t1597 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1976 VSS.t1578 a_867_n4378.t6 a_867_n7825.t1 VSS.t1575 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1977 VSS.t418 a_7272_2662.t4 a_7642_2662.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1978 a_5917_3666.t0 RWLB[0].t8 a_5465_n953.t26 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1979 a_2519_n5338.t1 Iref1.t2 a_2578_n5293.t1 VSS.t2221 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1980 VSS.t2158 a_6697_4148.t5 a_7067_4148.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1981 a_7752_2406.t2 WWL[5].t10 a_8020_4887.t2 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1982 a_8422_4686.t2 a_8327_4671.t3 VDD.t1503 VDD.t1502 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1983 a_7752_n286.t0 WWLD[4].t10 a_8020_4887.t16 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1984 a_4385_n1770.t2 a_4570_4887.t27 a_4578_n1770.t1 VSS.t227 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X1985 a_2683_n953.t13 WWL[4].t13 a_2672_2662.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1986 VSS.t1348 a_7847_693.t4 a_7752_678.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1987 VDD.t1045 a_n2415_n7216.t3 ADC1_OUT[2].t1 VDD.t1044 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1988 VSS.t1433 a_372_2662.t4 a_277_2647.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1989 VSS.t1172 a_2652_n2234.t3 a_2775_n2132.t0 VSS.t1171 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1990 a_7272_3666.t0 a_7177_3651.t4 VSS.t2345 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1991 a_1440_n953.t30 RWL[10].t8 a_1440_1216.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1992 a_7847_1216.t1 a_7752_1201.t4 VSS.t786 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1993 a_4877_678.t2 WWL[12].t11 a_5145_4887.t14 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1994 a_7067_3907.t0 VSS.t661 a_6615_n953.t6 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1995 VDD.t1882 a_8422_2943.t3 a_8327_2928.t1 VDD.t1881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1996 VSS.t890 a_7847_2421.t3 a_8217_2421.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1997 a_290_1939.t0 a_277_1924.t4 VSS.t457 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1998 a_1129_n7216.t0 PRE_CLSA.t54 VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X1999 a_852_3892.t2 WWLD[3].t11 a_1120_4887.t6 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2000 a_4192_1939.t0 RWLB[7].t6 a_3740_n953.t27 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2001 a_6615_4445.t1 a_6602_4430.t4 VSS.t1104 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2002 a_9367_2943.t1 RWLB[3].t3 a_8915_n953.t44 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2003 a_3152_2928.t0 WWL[3].t11 a_3420_4887.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2004 a_1522_n30.t0 a_1427_n45.t3 VSS.t1450 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2005 a_3258_n953.t1 WWL[5].t11 a_3247_2421.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2006 a_277_2165.t0 WWL[6].t12 a_545_4887.t19 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2007 VDD.t2238 a_7272_2180.t3 a_7177_2165.t1 VDD.t2237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2008 a_7847_4445.t1 a_7752_4430.t3 VDD.t1087 VDD.t1086 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2009 a_8422_1939.t1 a_8327_1924.t4 VSS.t2238 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2010 a_947_211.t0 a_852_196.t3 VSS.t463 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2011 a_12736_n5293.t1 VCLP.t44 a_12701_n5092.t0 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2012 a_4890_n953.t26 RWL[11].t3 a_4890_975.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2013 a_6040_n953.t15 VSS.t660 a_6040_n1053.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2014 a_947_1939.t1 a_852_1924.t4 VSS.t433 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2015 a_3701_n5338.t0 VCLP.t45 a_3563_n5338.t1 VSS.t203 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2016 VSS.t1390 a_947_3907.t3 a_1317_3907.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2017 a_4192_975.t0 RWLB[11].t7 a_3740_n953.t42 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2018 VSS.t311 SAEN.t34 a_902_n6503.t0 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2019 a_6492_3666.t0 RWLB[0].t9 a_6040_n953.t25 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2020 VSS.t470 a_372_2180.t4 a_742_2180.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2021 VSS.t1378 a_2097_n1053.t3 a_2467_n1053.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2022 a_3740_n953.t17 VSS.t659 a_3740_n512.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2023 a_4397_4445.t1 a_4302_4430.t5 VSS.t2484 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2024 a_5558_n953.t23 WWLD[2].t13 a_5547_4148.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2025 a_8433_n953.t1 WWL[2].t10 a_8422_3184.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2026 a_5465_452.t0 a_5452_437.t4 VSS.t1162 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2027 VDD.t792 a_3822_211.t3 a_3727_196.t0 VDD.t791 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2028 a_6065_n5338.t0 VCLP.t46 a_5927_n5338.t1 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2029 a_7765_n953.t31 RWL[0].t11 a_7765_3666.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2030 a_8217_693.t1 RWLB[12].t4 a_7765_n953.t20 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2031 a_383_n953.t16 WWL[13].t14 a_372_452.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2032 VSS.t994 a_1522_975.t4 a_1427_960.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2033 a_372_n1053.t0 a_277_n1068.t4 VSS.t1191 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2034 a_958_n953.t25 WWL[2].t11 a_947_3184.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2035 VDD.t1562 a_6697_1939.t3 a_6602_1924.t1 VDD.t1561 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2036 a_4315_3184.t1 a_4302_3169.t4 VSS.t1320 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2037 a_7642_1939.t1 RWLB[7].t7 a_7190_n953.t34 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2038 a_4448_n3770.t2 a_4675_n4483.t3 ADC7_OUT[0].t1 VSS.t1224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2039 a_2015_n953.t13 VSS.t658 a_2015_4686.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2040 a_7067_3425.t1 RWLB[1].t3 a_6615_n953.t33 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2041 VSS.t1825 a_1522_1698.t4 a_1892_1698.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2042 a_6708_n953.t1 WWL[5].t12 a_6697_2421.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2043 a_1427_1924.t2 WWL[7].t12 a_1695_4887.t18 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2044 a_2002_1442.t0 WWL[9].t14 a_2270_4887.t16 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2045 a_n3495_n8071.t0 SAEN.t35 a_n3298_n8026.t0 VSS.t312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2046 a_2672_4148.t1 a_2577_4133.t3 VDD.t1265 VDD.t1264 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2047 a_852_3410.t0 WWL[1].t12 a_1120_4887.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2048 a_5547_3184.t2 a_5452_3169.t3 VDD.t2102 VDD.t2101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2049 a_290_n953.t44 RWL[12].t7 a_290_693.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2050 a_7190_4445.t1 a_7177_4430.t4 VSS.t1862 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2051 VSS.t1587 a_4397_3666.t5 a_4302_3651.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2052 a_9008_n953.t10 WWL[3].t12 a_8997_2943.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2053 a_6040_n953.t18 RWL[9].t4 a_6040_1457.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2054 a_4408_n953.t24 WWL[13].t15 a_4397_452.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2055 VSS.t1567 a_947_n271.t3 a_1317_n271.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2056 VSS.t1462 a_1522_n812.t4 a_1892_n812.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2057 a_1028_n2086.t0 WE.t14 a_958_n953.t7 VSS.t2387 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2058 VDD.t2240 a_8997_n30.t4 a_8902_n45.t1 VDD.t2239 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2059 VDD.t1835 a_11776_n8583.t3 ADC13_OUT[3].t1 VDD.t1834 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2060 a_5857_n5850.t1 ADC8_OUT[1].t4 a_5927_n5338.t2 VSS.t1444 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2061 VSS.t314 SAEN.t36 a_10362_n3770.t0 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2062 a_2097_n812.t1 a_2002_n827.t3 VDD.t948 VDD.t947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2063 VSS.t1803 a_947_3425.t3 a_1317_3425.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2064 a_3822_2421.t0 a_3727_2406.t3 VDD.t562 VDD.t561 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2065 VSS.t1679 a_2097_1457.t3 a_2467_1457.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2066 a_2311_n7216.t2 ADC5_OUT[2].t4 a_2381_n7203.t2 VSS.t1103 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2067 VDD.t1833 SA_OUT[15].t3 a_8935_n1371.t1 VDD.t1832 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2068 VSS.t1996 a_5547_n1053.t3 a_5917_n1053.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2069 a_2097_3184.t1 a_2002_3169.t5 VSS.t2266 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2070 a_4315_n953.t39 RWL[12].t8 a_4315_693.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2071 a_1440_n953.t14 VSS.t657 a_1440_4445.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2072 a_7847_4445.t0 a_7752_4430.t4 VSS.t1374 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2073 a_3822_n271.t2 a_3727_n286.t3 VDD.t1015 VDD.t1014 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2074 VDD.t536 a_7847_2421.t4 a_7752_2406.t0 VDD.t535 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2075 VSS.t1220 a_3247_693.t4 a_3152_678.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2076 a_n1233_n8583.t1 ADC2_OUT[3].t3 VDD.t1640 VDD.t1639 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2077 a_n3565_n4483.t1 ADC0_OUT[0].t3 a_n3495_n4470.t2 VSS.t1164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2078 a_2097_693.t0 a_2002_678.t4 VSS.t1885 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2079 a_6040_n953.t48 RWL[14].t6 a_6040_211.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2080 a_5547_975.t2 a_5452_960.t4 VDD.t1077 VDD.t1076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2081 VDD.t1405 a_372_2421.t3 a_277_2406.t1 VDD.t1404 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2082 a_13864_n7216.t2 ADC15_OUT[2].t3 VDD.t1088 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2083 a_12963_n8583.t2 ADC14_OUT[3].t4 a_13033_n8071.t2 VSS.t1540 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2084 a_2590_2662.t1 a_2577_2647.t4 VSS.t1874 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 a_4972_2662.t0 a_4877_2647.t4 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2086 VSS.t1620 a_4972_211.t4 a_4877_196.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2087 VDD.t53 a_5547_211.t4 a_5452_196.t1 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2088 a_4877_3892.t2 WWLD[3].t12 a_5145_4887.t4 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2089 a_5452_1442.t0 WWL[9].t15 a_5720_4887.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2090 a_742_1457.t1 RWLB[9].t4 a_290_n953.t30 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2091 a_10589_n8583.t0 PRE_CLSA.t55 VDD.t197 VDD.t196 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2092 a_6812_n3770.t2 VCLP.t47 a_6777_n4116.t0 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2093 VSS.t1552 a_1522_1216.t4 a_1892_1216.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2094 a_7177_2928.t0 WWL[3].t13 a_7445_4887.t9 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2095 a_7283_n953.t2 WWL[5].t13 a_7272_2421.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2096 VDD.t515 a_947_3907.t4 a_852_3892.t0 VDD.t514 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2097 a_277_n45.t1 WWL[15].t14 a_545_4887.t16 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2098 a_7765_n953.t1 RWL[15].t4 a_7765_n30.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2099 a_947_n512.t2 a_852_n527.t3 VDD.t1402 VDD.t1401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2100 VSS.t1748 a_4972_3907.t4 a_5342_3907.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2101 a_3165_2421.t1 a_3152_2406.t5 VSS.t1838 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2102 VSS.t1812 a_5547_1457.t3 a_5917_1457.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2103 a_5547_3184.t1 a_5452_3169.t4 VSS.t2280 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2104 VSS.t1883 a_2672_975.t4 a_3042_975.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2105 VDD.t1011 a_2097_n1053.t4 a_2002_n1068.t0 VDD.t1010 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2106 a_3165_n271.t1 a_3152_n286.t5 VSS.t1877 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2107 a_2311_n5850.t0 PRE_CLSA.t56 VDD.t199 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2108 VSS.t1868 a_8997_3907.t5 a_8902_3892.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2109 a_4883_n5338.t1 Iref1.t3 a_4942_n5293.t1 VSS.t2222 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2110 VSS.t1863 a_6122_n1053.t4 a_6492_n1053.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2111 a_8433_n953.t22 WWL[15].t15 a_8422_n30.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2112 a_9405_n5850.t1 ADC11_OUT[1].t3 VDD.t1430 VDD.t1429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2113 a_1502_n2234.t0 Din[2].t1 VSS.t1760 VSS.t1759 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2114 a_3617_693.t1 RWLB[12].t5 a_3165_n953.t18 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2115 a_8902_n1068.t2 WWLD[7].t11 a_9170_4887.t25 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2116 VDD.t2187 a_3822_3666.t5 a_3727_3651.t1 VDD.t2186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2117 a_2002_4671.t2 WWLD[0].t14 a_2270_4887.t23 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2118 a_5465_4148.t1 a_5452_4133.t5 VSS.t934 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2119 a_8422_2662.t1 a_8327_2647.t3 VDD.t1695 VDD.t1694 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2120 VSS.t1077 a_6697_1698.t5 a_7067_1698.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2121 VSS.t1843 a_7272_n30.t3 a_7642_n30.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2122 a_7247_n5338.t1 Iref1.t4 a_7306_n5293.t1 VSS.t2223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2123 a_8327_3892.t2 WWLD[3].t13 a_8595_4887.t4 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2124 a_8340_3184.t0 a_8327_3169.t5 VSS.t382 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2125 a_7847_n30.t2 a_7752_n45.t3 VSS.t1796 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2126 a_6040_n953.t11 VSS.t656 a_6040_4686.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2127 a_5342_211.t1 RWLB[14].t7 a_4890_n953.t46 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2128 a_865_3184.t0 a_852_3169.t5 VSS.t1075 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2129 VDD.t1322 a_947_n271.t4 a_852_n286.t1 VDD.t1321 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2130 a_4877_3410.t0 WWL[1].t13 a_5145_4887.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2131 VSS.t1035 a_6697_n812.t5 a_7067_n812.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2132 a_11846_n8071.t0 SAEN.t37 a_12043_n8026.t0 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2133 a_4397_n512.t1 a_4302_n527.t3 VDD.t1346 VDD.t1345 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2134 VSS.t1200 a_8422_3666.t4 a_8327_3651.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2135 a_4767_3184.t1 RWLB[2].t10 a_4315_n953.t42 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2136 VSS.t1762 a_5527_n2234.t3 a_5650_n2132.t0 VSS.t1761 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2137 VSS.t839 a_2097_4686.t3 a_2467_4686.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2138 a_383_n953.t14 WWL[7].t13 a_372_1939.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2139 VSS.t971 a_4972_n271.t4 a_5342_n271.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2140 VSS.t2437 a_n1495_n4378.t5 a_n1495_n6849.t1 VSS.t2436 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2141 VDD.t1556 a_947_3425.t4 a_852_3410.t1 VDD.t1555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2142 a_6615_2421.t0 a_6602_2406.t4 VSS.t1418 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2143 VDD.t1418 a_2097_1457.t4 a_2002_1442.t1 VDD.t1417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2144 a_11549_n8026.t1 VCLP.t48 a_11514_n7825.t0 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2145 VDD.t1760 a_5547_n1053.t4 a_5452_n1068.t1 VDD.t1759 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2146 a_3822_2180.t1 a_3727_2165.t4 VSS.t989 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2147 VSS.t317 SAEN.t38 a_902_n3770.t0 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2148 a_4377_n2234.t1 Din[7].t1 VSS.t2016 VSS.t2015 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2149 VSS.t251 a_3822_693.t4 a_4192_693.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2150 a_8340_n30.t1 a_8327_n45.t5 VSS.t247 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2151 a_6615_n271.t1 a_6602_n286.t4 VSS.t113 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2152 VSS.t1611 a_8997_n271.t5 a_8902_n286.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2153 VSS.t1305 a_4972_3425.t4 a_5342_3425.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2154 VSS.t965 a_6122_1457.t4 a_6492_1457.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2155 VDD.t77 a_n52_n8583.t3 ADC3_OUT[3].t2 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2156 a_3833_n953.t9 WWLD[3].t14 a_3822_3907.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2157 a_7847_2421.t2 a_7752_2406.t3 VDD.t1884 VDD.t1883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2158 VDD.t566 a_12963_n5850.t3 ADC14_OUT[1].t1 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2159 a_1317_n812.t0 VSS.t655 a_865_n953.t14 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2160 a_1120_4887.t25 PRE_SRAM.t19 VDD.t2045 VDD.t2044 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2161 a_1533_n953.t4 WWL[11].t13 a_1522_975.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2162 a_4972_452.t1 a_4877_437.t4 VDD.t1300 VDD.t1299 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2163 a_7847_n271.t2 a_7752_n286.t3 VDD.t2263 VDD.t2262 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2164 a_1199_n8071.t0 SAEN.t39 a_1396_n8026.t0 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2165 VDD.t201 PRE_CLSA.t57 ADC6_OUT[3].t0 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2166 VSS.t1089 a_8997_3425.t5 a_8902_3410.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2167 VSS.t2316 a_7843_n2422.t5 a_11514_n6849.t0 VSS.t2315 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2168 a_156_n8071.t1 Iref3.t10 a_215_n8026.t1 VSS.t829 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2169 a_4983_n953.t20 WWLD[7].t12 a_4972_n1053.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2170 a_5452_4671.t2 WWLD[0].t15 a_5720_4887.t5 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2171 a_8915_4148.t1 a_8902_4133.t3 VSS.t1403 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2172 a_1440_n953.t48 RWL[14].t7 a_1440_211.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2173 VSS.t1009 a_8402_n2234.t3 a_8525_n2132.t0 VSS.t1008 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2174 a_742_4686.t0 VSS.t654 a_290_n953.t6 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2175 a_8997_2180.t1 a_8902_2165.t5 VDD.t1618 VDD.t1617 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 VSS.t1522 a_1522_4445.t4 a_1892_4445.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2177 a_9008_n953.t13 WWL[15].t16 a_8997_n30.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2178 a_2652_n2234.t1 Din[4].t1 VSS.t1283 VSS.t1282 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2179 a_4397_2421.t1 a_4302_2406.t5 VSS.t1095 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2180 VSS.t1030 a_6697_1216.t5 a_7067_1216.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2181 a_4408_n953.t20 WWL[0].t11 a_4397_3666.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2182 a_8327_3410.t0 WWL[1].t14 a_8595_4887.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2183 a_5558_n953.t5 WWL[8].t13 a_5547_1698.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 a_4397_n271.t0 a_4302_n286.t5 VSS.t1085 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2185 VSS.t987 a_6693_n2422.t6 a_9143_n7825.t1 VSS.t984 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2186 a_7039_n4483.t0 PRE_CLSA.t58 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2187 VSS.t1644 a_7847_n30.t4 a_8217_n30.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2188 VSS.t414 a_5547_4686.t3 a_5917_4686.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2189 VDD.t343 a_8422_3907.t3 a_8327_3892.t0 VDD.t342 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2190 VDD.t1566 a_5547_1457.t4 a_5452_1442.t2 VDD.t1565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2191 a_3740_n953.t5 RWL[15].t5 a_3740_n30.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2192 a_2015_n953.t45 RWL[4].t4 a_2015_2662.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2193 VDD.t1988 a_6122_975.t3 a_6027_960.t1 VDD.t1987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2194 a_5558_n953.t17 WWLD[6].t18 a_5547_n812.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2195 a_2381_n5338.t0 SAEN.t40 a_2578_n5293.t0 VSS.t291 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2196 a_2311_n4483.t1 ADC5_OUT[0].t3 a_2381_n4470.t2 VSS.t1126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2197 a_7190_2421.t1 a_7177_2406.t5 VSS.t2377 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2198 VDD.t2191 a_947_452.t5 a_852_437.t1 VDD.t2190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2199 a_3833_n953.t15 WWLD[4].t11 a_3822_n271.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2200 a_13864_n7216.t0 PRE_CLSA.t59 VDD.t204 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2201 a_6697_4148.t0 a_6602_4133.t5 VSS.t1097 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2202 a_1522_3666.t1 a_1427_3651.t3 VDD.t904 VDD.t903 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2203 a_2672_1698.t1 a_2577_1683.t3 VDD.t1861 VDD.t1860 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2204 a_6697_211.t2 a_6602_196.t3 VDD.t1008 VDD.t1007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2205 a_7190_n271.t1 a_7177_n286.t5 VSS.t2352 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2206 a_5527_n2234.t1 Din[9].t1 VSS.t2103 VSS.t2102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2207 VDD.t730 a_4972_n512.t3 a_4877_n527.t0 VDD.t729 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2208 a_4983_n953.t21 WWL[9].t16 a_4972_1457.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2209 a_6602_678.t2 WWL[12].t12 a_6870_4887.t10 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2210 a_3833_n953.t2 WWL[1].t15 a_3822_3425.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2211 a_10589_n5850.t1 ADC12_OUT[1].t4 a_10659_n5338.t2 VSS.t1542 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2212 a_3903_n2086.t0 WE.t15 a_3833_n953.t14 VSS.t2388 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2213 VSS.t1740 a_8997_n512.t3 a_9367_n512.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2214 a_6122_n812.t1 a_6027_n827.t4 VSS.t886 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2215 a_1440_n953.t47 RWL[5].t9 a_1440_2421.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2216 a_7847_2421.t1 a_7752_2406.t4 VSS.t2128 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2217 a_7039_n7216.t2 ADC9_OUT[2].t4 a_7109_n7203.t2 VSS.t1939 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2218 a_7847_n271.t1 a_7752_n286.t4 VSS.t2496 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2219 a_2519_n7203.t1 Iref2.t2 a_2578_n6847.t1 VSS.t1980 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2220 a_2590_2943.t1 a_2577_2928.t5 VSS.t2242 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2221 VDD.t646 a_8422_n271.t3 a_8327_n286.t0 VDD.t645 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2222 VDD.t496 a_2097_4686.t4 a_2002_4671.t0 VDD.t495 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2223 a_4972_2943.t2 a_4877_2928.t4 VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2224 a_2015_n30.t1 a_2002_n45.t4 VSS.t1362 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2225 a_2127_n1770.t0 a_2108_n953.t27 a_2085_n1770.t1 VSS.t2153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2226 a_5558_n953.t7 WWL[10].t14 a_5547_1216.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2227 VSS.t1492 a_5632_n6430# a_9178_n6503.t0 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2228 a_6102_n2234.t0 Din[10].t0 VDD.t1006 VDD.t1005 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2229 a_8792_3184.t1 RWLB[2].t11 a_8340_n953.t44 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 a_3617_n512.t0 VSS.t653 a_3165_n953.t6 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2231 VSS.t2111 a_6122_4686.t4 a_6492_4686.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2232 VDD.t630 a_8422_3425.t3 a_8327_3410.t1 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2233 a_2577_3169.t0 WWL[2].t12 a_2845_4887.t24 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2234 VDD.t998 a_5857_n8583.t3 ADC8_OUT[3].t1 VDD.t997 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2235 a_4890_n953.t38 RWL[6].t4 a_4890_2180.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2236 a_3740_n953.t8 VSS.t652 a_3740_4148.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2237 a_9008_n953.t3 WWLD[3].t15 a_8997_3907.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2238 a_6778_n2086.t1 WE.t16 a_6708_n953.t6 VSS.t2389 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2239 a_3740_n30.t1 a_3727_n45.t5 VSS.t2212 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2240 a_4315_n953.t2 RWL[15].t6 a_4315_n30.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2241 a_8595_4887.t22 PRE_SRAM.t20 VDD.t2047 VDD.t2046 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2242 a_2672_1216.t0 a_2577_1201.t3 VDD.t654 VDD.t653 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2243 VDD.t700 a_8221_n8583.t3 ADC10_OUT[3].t2 VDD.t699 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2244 a_5342_n812.t0 VSS.t651 a_4890_n953.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2245 VSS.t1712 a_6697_4445.t5 a_7067_4445.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2246 a_3740_3907.t1 a_3727_3892.t5 VSS.t2262 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2247 a_2015_1939.t0 a_2002_1924.t4 VSS.t1707 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 a_n1163_n7203.t0 SAEN.t41 a_n966_n6847.t0 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2249 a_6122_3907.t1 a_6027_3892.t3 VDD.t982 VDD.t981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2250 VSS.t1559 a_6697_3184.t4 a_6602_3169.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2251 VSS.t2156 a_1522_2180.t4 a_1427_2165.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2252 a_5465_n953.t29 RWL[7].t9 a_5465_1939.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2253 a_7858_n953.t4 WWLD[5].t19 a_7847_n512.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2254 a_8217_2180.t0 RWLB[6].t5 a_7765_n953.t26 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2255 a_3247_1939.t1 a_3152_1924.t3 VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2256 a_8327_678.t1 WWL[12].t13 a_8595_4887.t5 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2257 VSS.t319 SAEN.t42 a_n2642_n6503.t0 VSS.t302 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2258 VDD.t345 a_5547_4686.t4 a_5452_4671.t0 VDD.t344 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2259 a_8422_2943.t2 a_8327_2928.t3 VDD.t1855 VDD.t1854 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2260 a_8433_n953.t26 WWL[0].t12 a_8422_3666.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2261 a_1695_4887.t5 PRE_SRAM.t21 a_1533_n953.t6 VDD.t2048 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2262 a_3266_n8026.t2 a_3493_n8583.t4 ADC6_OUT[3].t1 VSS.t1376 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2263 a_958_n953.t17 WWL[0].t13 a_947_3666.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2264 VSS.t1002 a_3247_2943.t3 a_3617_2943.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2265 a_2002_2647.t2 WWL[4].t14 a_2270_4887.t17 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2266 a_290_n512.t1 a_277_n527.t5 VSS.t2264 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2267 a_n2415_n7216.t0 PRE_CLSA.t60 VDD.t205 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2268 a_4315_3666.t1 a_4302_3651.t4 VSS.t2057 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2269 a_6040_n953.t45 RWL[4].t5 a_6040_2662.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2270 a_5465_1698.t1 a_5452_1683.t5 VSS.t1483 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2271 a_9008_n953.t19 WWLD[4].t12 a_8997_n271.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2272 a_4192_n512.t0 VSS.t650 a_3740_n953.t13 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2273 VSS.t2040 a_2097_1939.t5 a_2002_1924.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2274 a_7252_n2234.t1 Din[12].t0 VDD.t1434 VDD.t1433 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2275 a_360_n1770.t2 a_545_4887.t27 a_553_n1770.t1 VSS.t2306 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2276 a_4983_n953.t7 WWLD[0].t16 a_4972_4686.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2277 a_5547_3666.t1 a_5452_3651.t3 VDD.t966 VDD.t965 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2278 a_9008_n953.t0 WWL[1].t16 a_8997_3425.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2279 a_7642_975.t1 RWLB[11].t8 a_7190_n953.t41 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 a_8422_n512.t1 a_8327_n527.t4 VSS.t2154 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2281 VSS.t1512 a_2097_2662.t3 a_2467_2662.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2282 a_2002_196.t0 WWL[14].t15 a_2270_4887.t12 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2283 a_7928_n2086.t0 WE.t17 a_7858_n953.t8 VSS.t2390 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2284 VDD.t1485 a_8997_n512.t4 a_8902_n527.t2 VDD.t1484 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2285 a_7765_n953.t25 RWL[14].t8 a_7765_211.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 a_947_n512.t1 a_852_n527.t4 VSS.t1677 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2287 a_3563_n8071.t0 SAEN.t43 a_3760_n8026.t0 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2288 VSS.t321 SAEN.t44 a_12736_n5293.t0 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2289 a_8915_n953.t32 RWL[7].t10 a_8915_1939.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2290 a_8915_452.t0 a_8902_437.t4 VSS.t841 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2291 VSS.t1739 a_6697_211.t3 a_6602_196.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2292 VDD.t2050 PRE_SRAM.t22 a_2683_n953.t22 VDD.t2049 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2293 a_2097_3666.t0 a_2002_3651.t5 VSS.t1795 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2294 a_3740_3425.t0 a_3727_3410.t5 VSS.t2498 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2295 a_6697_1939.t2 a_6602_1924.t3 VDD.t1013 VDD.t1012 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2296 a_4890_1457.t0 a_4877_1442.t5 VSS.t2210 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2297 a_5558_n953.t24 WWLD[1].t14 a_5547_4445.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2298 a_6122_3425.t2 a_6027_3410.t3 VDD.t1843 VDD.t1842 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2299 a_7272_1457.t0 a_7177_1442.t3 VDD.t438 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2300 a_2097_452.t0 a_2002_437.t3 VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2301 a_5927_n8071.t0 SAEN.t45 a_6124_n8026.t0 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2302 a_5452_2647.t2 WWL[4].t15 a_5720_4887.t19 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2303 VDD.t207 PRE_CLSA.t61 ADC10_OUT[3].t0 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2304 a_290_n953.t42 RWL[3].t4 a_290_2943.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2305 a_902_n5293.t2 a_1129_n5850.t4 ADC4_OUT[1].t2 VSS.t1521 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2306 a_7752_3169.t2 WWL[2].t13 a_8020_4887.t23 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2307 a_742_2662.t1 RWLB[4].t4 a_290_n953.t37 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2308 VSS.t1681 a_1522_2421.t4 a_1892_2421.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2309 a_8915_1698.t0 a_8902_1683.t3 VSS.t416 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2310 VSS.t2007 a_3822_2943.t3 a_4192_2943.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2311 VSS.t1683 a_5547_1939.t5 a_5452_1924.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2312 VDD.t1942 a_7272_452.t4 a_7177_437.t2 VDD.t1941 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2313 a_5630_n8026.t1 VCLP.t49 a_5595_n7825.t0 VSS.t207 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2314 a_7642_n512.t0 VSS.t649 a_7190_n953.t13 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2315 a_4972_3907.t0 a_4877_3892.t3 VSS.t770 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2316 a_3247_1939.t0 a_3152_1924.t4 VSS.t439 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2317 a_1427_n527.t0 WWLD[5].t20 a_1695_4887.t14 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2318 a_2672_4445.t1 a_2577_4430.t3 VDD.t1436 VDD.t1435 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2319 a_5465_1216.t1 a_5452_1201.t5 VSS.t1562 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2320 a_n3565_n7216.t0 PRE_CLSA.t62 VDD.t208 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2321 VSS.t1124 a_5547_2662.t3 a_5917_2662.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2322 a_4745_n5338.t0 SAEN.t46 a_4942_n5293.t0 VSS.t296 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2323 VSS.t1020 a_n2677_n4378.t0 a_n2677_n4378.t1 VSS.t1019 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2324 VSS.t1001 a_7847_3184.t3 a_8217_3184.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2325 VSS.t2082 a_2672_2180.t4 a_3042_2180.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 VSS.t1829 a_8422_452.t4 a_8327_437.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2327 VSS.t783 a_5118_n2426.t5 a_5595_n6849.t0 VSS.t782 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2328 a_3258_n953.t15 WWL[12].t14 a_3247_693.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2329 a_7190_n1053.t1 a_7177_n1068.t4 VSS.t1904 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2330 a_6602_n827.t0 WWLD[6].t19 a_6870_4887.t19 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2331 a_5002_n1770.t0 SA_OUT[8].t4 a_4910_n1371.t0 VSS.t1659 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2332 VDD.t1711 SA_OUT[1].t3 a_885_n1371.t1 VDD.t1710 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2333 a_3258_n953.t24 WWL[2].t14 a_3247_3184.t1 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2334 a_6040_1939.t1 a_6027_1924.t5 VSS.t977 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2335 a_7109_n5338.t0 SAEN.t47 a_7306_n5293.t0 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2336 a_n1025_n5338.t0 VCLP.t50 a_n1163_n5338.t1 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2337 a_7039_n4483.t1 ADC9_OUT[0].t3 a_7109_n4470.t2 VSS.t1504 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2338 a_5547_3666.t0 a_5452_3651.t4 VSS.t1325 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2339 a_6697_1698.t1 a_6602_1683.t5 VSS.t1000 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2340 a_156_n5338.t0 VCLP.t51 a_18_n5338.t1 VSS.t209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2341 a_3727_196.t1 WWL[14].t16 a_3995_4887.t19 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2342 VDD.t210 PRE_CLSA.t63 ADC15_OUT[3].t0 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2343 VDD.t212 PRE_CLSA.t64 ADC3_OUT[1].t0 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2344 VDD.t494 a_1522_1939.t3 a_1427_1924.t0 VDD.t493 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2345 a_5547_693.t2 a_5452_678.t3 VSS.t2278 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2346 VDD.t628 a_3247_2943.t4 a_3152_2928.t1 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2347 a_4983_n953.t10 WWL[12].t15 a_4972_693.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2348 a_6027_2165.t2 WWL[6].t13 a_6295_4887.t25 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2349 a_2467_1939.t1 RWLB[7].t8 a_2015_n953.t35 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2350 a_8902_960.t0 WWL[11].t14 a_9170_4887.t26 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2351 a_4883_n7203.t1 Iref2.t3 a_4942_n6847.t1 VSS.t1981 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2352 VSS.t324 SAEN.t48 a_9178_n3770.t0 VSS.t323 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2353 VSS.t1735 a_7272_2943.t4 a_7642_2943.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2354 a_7272_211.t2 a_7177_196.t3 VSS.t2488 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2355 a_1317_975.t0 RWLB[11].t9 a_865_n953.t41 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2356 a_n2415_n8583.t2 ADC1_OUT[3].t4 a_n2345_n8071.t2 VSS.t1661 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2357 a_5465_n1053.t0 a_5452_n1068.t4 VSS.t767 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2358 a_8340_3666.t0 a_8327_3651.t5 VSS.t1272 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2359 a_8915_1216.t1 a_8902_1201.t3 VSS.t2014 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2360 a_7067_452.t0 RWLB[13].t7 a_6615_n953.t20 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2361 a_3277_n1770.t1 SA_OUT[5].t4 a_3185_n1371.t1 VSS.t408 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2362 VSS.t2065 a_6122_1939.t4 a_6027_1924.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2363 a_4315_n953.t17 VSS.t648 a_4315_n1053.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2364 VDD.t1262 a_2097_2662.t4 a_2002_2647.t0 VDD.t1261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2365 a_6040_693.t1 a_6027_678.t5 VSS.t975 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2366 a_7247_n7203.t1 Iref2.t4 a_7306_n6847.t1 VSS.t1982 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2367 a_865_3666.t0 a_852_3651.t5 VSS.t1392 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2368 a_4972_3425.t1 a_4877_3410.t3 VSS.t1303 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2369 a_2683_n953.t11 WWL[3].t14 a_2672_2943.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2370 a_3247_n30.t2 a_3152_n45.t4 VDD.t1734 VDD.t1733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2371 VSS.t1136 a_372_2943.t4 a_277_2928.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2372 a_5002_n1770.t1 a_4983_n953.t27 a_4960_n1770.t0 VSS.t2118 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2373 VSS.t1744 a_6122_2662.t4 a_6492_2662.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2374 a_4767_3666.t0 RWLB[0].t10 a_4315_n953.t24 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2375 a_8792_452.t0 RWLB[13].t8 a_8340_n953.t24 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2376 VDD.t1316 a_10589_n8583.t3 ADC12_OUT[3].t1 VDD.t1315 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2377 a_n1163_n4470.t0 SAEN.t49 a_n966_n4114.t0 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2378 a_4890_4686.t1 a_4877_4671.t5 VSS.t2287 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2379 a_6708_n953.t25 WWL[2].t15 a_6697_3184.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2380 a_1533_n953.t11 WWL[6].t14 a_1522_2180.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2381 a_7272_4686.t1 a_7177_4671.t3 VDD.t1244 VDD.t1243 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2382 a_3740_n953.t31 RWL[8].t7 a_3740_1698.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2383 VSS.t327 SAEN.t50 a_n2642_n3770.t0 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2384 VSS.t1964 a_947_n1053.t5 a_852_n1068.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2385 a_8340_n1053.t1 a_8327_n1068.t4 VSS.t964 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2386 a_6697_1216.t0 a_6602_1201.t5 VSS.t1775 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2387 a_6152_n1770.t0 SA_OUT[10].t4 a_6060_n1371.t1 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2388 VDD.t753 SA_OUT[3].t3 a_2035_n1371.t0 VDD.t752 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2389 a_5917_1939.t0 RWLB[7].t9 a_5465_n953.t38 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2390 a_3740_n953.t14 VSS.t647 a_3740_n812.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2391 VSS.t1800 a_6697_2421.t5 a_7067_2421.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2392 a_3042_1457.t0 RWLB[9].t5 a_2590_n953.t29 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2393 a_3165_n953.t42 RWL[13].t5 a_3165_452.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2394 a_8902_4133.t0 WWLD[2].t14 a_9170_4887.t13 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2395 a_3822_3184.t1 a_3727_3169.t3 VDD.t890 VDD.t889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2396 a_2108_n953.t14 WWL[7].t14 a_2097_1939.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2397 a_9613_n8071.t1 Iref3.t11 a_9672_n8026.t1 VSS.t830 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2398 a_7877_n1770.t1 a_7858_n953.t27 a_7835_n1770.t2 VSS.t2301 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2399 a_5465_4445.t1 a_5452_4430.t5 VSS.t899 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2400 a_4315_n953.t19 RWL[9].t5 a_4315_1457.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2401 a_2002_2928.t0 WWL[3].t15 a_2270_4887.t14 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2402 VDD.t745 a_5547_2662.t4 a_5452_2647.t0 VDD.t744 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2403 VSS.t1472 a_2097_452.t4 a_2002_437.t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2404 VDD.t442 a_2672_452.t4 a_2577_437.t0 VDD.t441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2405 VDD.t1720 a_6122_2180.t3 a_6027_2165.t0 VDD.t1719 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2406 a_7272_1939.t1 a_7177_1924.t4 VSS.t1455 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2407 VDD.t1718 a_4972_4148.t3 a_4877_4133.t2 VDD.t1717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2408 VDD.t339 a_7847_3184.t4 a_7752_3169.t0 VDD.t338 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2409 a_6615_n1053.t1 a_6602_n1068.t3 VSS.t1909 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 VDD.t1438 a_372_3184.t3 a_277_3169.t2 VDD.t1437 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2411 a_4890_n953.t47 RWL[13].t6 a_4890_452.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2412 a_4427_n1770.t0 SA_OUT[7].t4 a_4335_n1371.t0 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2413 VSS.t2025 a_8997_4148.t3 a_9367_4148.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2414 VSS.t1733 a_7272_693.t3 a_7642_693.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2415 a_1129_n8583.t2 ADC4_OUT[3].t4 a_1199_n8071.t2 VSS.t1046 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2416 VSS.t1066 a_3231_n4378.t5 a_3231_n4116.t1 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2417 a_4983_n953.t22 WWL[4].t16 a_4972_2662.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2418 VSS.t1190 a_947_1457.t5 a_852_1442.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2419 a_2590_n953.t16 VSS.t646 a_2590_n512.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2420 a_8422_452.t1 a_8327_437.t4 VDD.t574 VDD.t573 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2421 a_7283_n953.t26 WWL[2].t16 a_7272_3184.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2422 a_3740_n953.t2 RWL[10].t9 a_3740_1216.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2423 a_9367_3907.t0 VSS.t645 a_8915_n953.t10 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2424 a_3152_3892.t2 WWLD[3].t16 a_3420_4887.t9 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2425 a_3165_3184.t0 a_3152_3169.t5 VSS.t1259 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2426 VSS.t1926 a_n314_n4378.t5 a_n314_n4116.t1 VSS.t1922 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2427 a_8915_4445.t1 a_8902_4430.t3 VSS.t2012 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2428 a_6492_1939.t0 RWLB[7].t10 a_6040_n953.t38 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2429 a_4302_960.t0 WWL[11].t15 a_4570_4887.t26 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2430 a_5452_2928.t2 WWL[3].t16 a_5720_4887.t16 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2431 a_5558_n953.t10 WWL[5].t14 a_5547_2421.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2432 a_2672_211.t0 a_2577_196.t3 VSS.t497 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2433 a_2002_n1068.t2 WWLD[7].t13 a_2270_4887.t15 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2434 a_742_2943.t0 RWLB[3].t4 a_290_n953.t34 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2435 a_2467_452.t1 RWLB[13].t9 a_2015_n953.t19 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2436 a_947_n30.t1 a_852_n45.t3 VSS.t1715 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2437 a_13637_n8026.t2 a_13864_n8583.t4 ADC15_OUT[3].t2 VSS.t1409 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2438 a_8340_n953.t19 VSS.t644 a_8340_n1053.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2439 VSS.t2370 a_3247_3907.t3 a_3617_3907.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2440 a_1440_693.t1 a_1427_678.t5 VSS.t422 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2441 a_372_1457.t1 a_277_1442.t4 VSS.t916 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2442 VSS.t797 a_947_975.t3 a_1317_975.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2443 a_n52_n7216.t0 PRE_CLSA.t65 VDD.t213 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2444 a_865_n953.t8 VSS.t643 a_865_n1053.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2445 a_10362_n8026.t1 VCLP.t52 a_10327_n7825.t0 VSS.t210 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2446 a_8792_3666.t0 RWLB[0].t11 a_8340_n953.t27 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2447 VSS.t2209 a_3822_n30.t4 a_4192_n30.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2448 a_947_n812.t2 a_852_n827.t3 VDD.t1634 VDD.t1633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2449 a_2672_2421.t0 a_2577_2406.t3 VDD.t578 VDD.t577 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2450 VSS.t2442 a_4397_n1053.t3 a_4767_n1053.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2451 a_7858_n953.t18 WWLD[2].t15 a_7847_4148.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2452 a_2577_3651.t2 WWL[0].t14 a_2845_4887.t25 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2453 VSS.t1157 a_6268_n2426.t5 a_7959_n6849.t0 VSS.t1156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2454 a_6697_4445.t0 a_6602_4430.t5 VSS.t1105 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2455 a_2672_n271.t0 a_2577_n286.t3 VDD.t826 VDD.t825 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2456 VDD.t1610 a_11776_n5850.t3 ADC13_OUT[1].t1 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2457 VSS.t2371 a_4972_n1053.t5 a_4877_n1068.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2458 a_3042_4686.t0 VSS.t642 a_2590_n953.t14 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2459 a_4877_n1068.t2 WWLD[7].t14 a_5145_4887.t25 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2460 a_1440_2180.t1 a_1427_2165.t5 VSS.t1640 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2461 VSS.t2133 a_7418_n2426.t5 a_10327_n6849.t0 VSS.t2132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2462 a_6615_3184.t1 a_6602_3169.t4 VSS.t1276 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2463 a_4315_n953.t11 VSS.t641 a_4315_4686.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2464 a_9367_3425.t0 RWLB[1].t4 a_8915_n953.t33 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2465 a_n1233_n5850.t1 ADC2_OUT[1].t3 VDD.t1776 VDD.t1775 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2466 a_3152_3410.t0 WWL[1].t17 a_3420_4887.t2 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2467 a_7847_3184.t2 a_7752_3169.t3 VDD.t474 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2468 a_4302_1442.t0 WWL[9].t17 a_4570_4887.t13 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2469 VSS.t2347 a_2672_n512.t4 a_2577_n527.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2470 a_6133_n953.t8 WWL[7].t15 a_6122_1939.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2471 VSS.t1933 a_6697_3666.t4 a_6602_3651.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2472 a_8340_n953.t22 RWL[9].t6 a_8340_1457.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2473 VSS.t1249 a_947_693.t3 a_1317_693.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2474 VSS.t2199 a_3247_n271.t3 a_3617_n271.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2475 a_9405_n5850.t2 ADC11_OUT[1].t4 a_9475_n5338.t1 VSS.t905 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2476 VSS.t2275 a_1502_n2234.t4 a_1625_n2132.t0 VSS.t2274 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2477 VDD.t1782 a_8997_4148.t4 a_8902_4133.t1 VDD.t1781 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2478 a_290_n953.t12 VSS.t640 a_290_3907.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2479 a_865_n953.t21 RWL[9].t7 a_865_1457.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2480 a_6027_960.t0 WWL[11].t16 a_6295_4887.t3 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2481 a_10589_n5850.t0 PRE_CLSA.t66 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2482 a_3152_n1068.t2 WWLD[7].t15 a_3420_4887.t20 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 VSS.t1301 a_2672_211.t5 a_3042_211.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2484 VSS.t1506 a_4397_n30.t4 a_4302_n45.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2485 VSS.t1117 a_947_4686.t5 a_852_4671.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2486 VSS.t2446 a_3822_3907.t3 a_4192_3907.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2487 VSS.t2451 a_3247_3425.t3 a_3617_3425.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2488 VSS.t1415 a_4397_1457.t3 a_4767_1457.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2489 a_4397_n812.t1 a_4302_n827.t3 VDD.t1930 VDD.t1929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2490 a_4397_3184.t1 a_4302_3169.t5 VSS.t1321 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2491 a_7994_n5293.t1 VCLP.t53 a_7959_n5092.t0 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2492 a_3740_n953.t12 VSS.t639 a_3740_4445.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2493 VSS.t2217 a_4972_1457.t5 a_4877_1442.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2494 a_3822_452.t2 a_3727_437.t4 VDD.t1103 VDD.t1102 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 VSS.t1208 a_5543_n2422.t2 a_5543_n2422.t3 VSS.t1207 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2496 a_4890_2662.t1 a_4877_2647.t5 VSS.t1692 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2497 a_7190_3184.t0 a_7177_3169.t5 VSS.t1466 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2498 a_7272_2662.t0 a_7177_2647.t3 VDD.t884 VDD.t883 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2499 a_3493_n7216.t0 ADC6_OUT[2].t4 a_3563_n7203.t1 VSS.t1424 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2500 a_7177_3892.t0 WWLD[3].t17 a_7445_4887.t4 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2501 a_8221_n8583.t0 ADC10_OUT[3].t3 VDD.t349 VDD.t348 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2502 a_6027_n1068.t2 WWLD[7].t16 a_6295_4887.t19 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2503 a_2015_n512.t1 a_2002_n527.t4 VSS.t1994 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2504 a_13934_n7203.t1 a_5632_n6430# a_14131_n6847.t0 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2505 a_12736_n5293.t2 a_12963_n5850.t4 ADC14_OUT[1].t2 VSS.t917 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2506 VDD.t2174 a_3247_3907.t4 a_3152_3892.t1 VDD.t2173 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2507 a_290_n953.t18 VSS.t638 a_290_n271.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2508 a_3247_n512.t0 a_3152_n527.t3 VDD.t315 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2509 a_372_4686.t0 a_277_4671.t4 VSS.t1527 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2510 VDD.t1293 a_947_975.t4 a_852_960.t2 VDD.t1292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2511 VSS.t1684 a_3822_n271.t3 a_4192_n271.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2512 VDD.t624 a_7039_n7216.t3 ADC9_OUT[2].t1 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2513 VSS.t2268 a_7272_3907.t4 a_7642_3907.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2514 a_5465_2421.t0 a_5452_2406.t5 VSS.t1133 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2515 VDD.t2213 a_4397_n1053.t4 a_4302_n1068.t2 VDD.t2212 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2516 a_1522_4148.t0 a_1427_4133.t4 VSS.t1844 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2517 a_7752_3651.t2 WWL[0].t15 a_8020_4887.t24 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2518 a_290_n953.t22 RWL[1].t4 a_290_3425.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2519 a_1440_n953.t24 RWL[2].t11 a_1440_3184.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2520 a_7847_3184.t1 a_7752_3169.t4 VSS.t805 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2521 a_2672_2180.t0 a_2577_2165.t4 VSS.t1524 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2522 a_8902_1683.t0 WWL[8].t14 a_9170_4887.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2523 VSS.t2000 a_4972_975.t4 a_5342_975.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2524 a_10797_n8071.t1 Iref3.t12 a_10856_n8026.t1 VSS.t831 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2525 a_5465_n271.t1 a_5452_n286.t5 VSS.t1144 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2526 VSS.t2494 a_3822_3425.t3 a_4192_3425.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2527 VSS.t1916 a_8422_n1053.t4 a_8792_n1053.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2528 a_2683_n953.t4 WWLD[3].t18 a_2672_3907.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2529 VSS.t1686 a_8997_975.t5 a_8902_960.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2530 VDD.t83 a_4972_1698.t4 a_4877_1683.t1 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2531 a_5452_196.t2 WWL[14].t17 a_5720_4887.t13 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2532 VSS.t2471 a_372_3907.t5 a_277_3892.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2533 VDD.t217 PRE_CLSA.t67 ADC13_OUT[3].t0 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2534 VDD.t878 a_n52_n5850.t3 ADC3_OUT[1].t1 VDD.t877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2535 VSS.t2141 a_8997_1698.t3 a_9367_1698.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2536 a_3493_n7216.t2 PRE_CLSA.t68 VDD.t218 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2537 a_4302_4671.t0 WWLD[0].t17 a_4570_4887.t18 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2538 a_7765_4148.t1 a_7752_4133.t5 VSS.t1339 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2539 VSS.t1849 a_7847_3666.t3 a_8217_3666.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2540 VDD.t37 a_4972_n812.t4 a_4877_n827.t1 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2541 VSS.t1932 a_7847_n512.t5 a_7752_n527.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2542 a_2015_n953.t46 RWL[3].t5 a_2015_2943.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2543 a_8997_211.t0 a_8902_196.t4 VSS.t2119 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2544 VDD.t220 PRE_CLSA.t69 ADC6_OUT[1].t0 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2545 VDD.t1788 SA_OUT[13].t3 a_7785_n1371.t1 VDD.t1787 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2546 a_8340_n953.t14 VSS.t637 a_8340_4686.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2547 a_5342_n30.t1 RWLB[15].t8 a_4890_n953.t43 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2548 VDD.t222 PRE_CLSA.t70 ADC14_OUT[0].t0 VDD.t221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2549 VDD.t2271 a_3227_n2234.t3 a_3350_n2132.t1 VDD.t2270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2550 VDD.t1129 PRE_VLSA.t25 a_885_n1371.t0 VDD.t1128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2551 a_372_2180.t0 a_277_2165.t3 VDD.t418 VDD.t417 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2552 VDD.t2223 a_3247_n271.t4 a_3152_n286.t1 VDD.t2222 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2553 VSS.t2208 a_8997_n812.t3 a_9367_n812.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2554 a_865_n953.t11 VSS.t636 a_865_4686.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2555 a_3258_n953.t25 WWL[0].t16 a_3247_3666.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2556 a_7177_3410.t0 WWL[1].t18 a_7445_4887.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2557 a_6697_n512.t1 a_6602_n527.t3 VDD.t2273 VDD.t2272 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2558 a_1892_2180.t0 RWLB[6].t6 a_1440_n953.t40 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2559 a_7765_693.t0 a_7752_678.t5 VSS.t1327 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2560 a_2077_n2234.t0 Din[3].t0 VDD.t1053 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2561 VSS.t2349 a_7272_n271.t4 a_7642_n271.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2562 VSS.t1012 a_4397_4686.t3 a_4767_4686.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2563 VDD.t2217 a_3247_3425.t4 a_3152_3410.t2 VDD.t2216 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2564 VDD.t1595 a_4397_1457.t4 a_4302_1442.t1 VDD.t1594 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2565 VDD.t1079 a_6697_n30.t5 a_6602_n45.t1 VDD.t1078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2566 a_9613_n5338.t0 VCLP.t54 a_9475_n5338.t2 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2567 a_8915_2421.t0 a_8902_2406.t3 VSS.t1420 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2568 a_3247_975.t1 a_3152_960.t3 VSS.t1288 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2569 a_947_693.t2 a_852_678.t4 VDD.t2236 VDD.t2235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2570 a_1427_960.t0 WWL[11].t17 a_1695_4887.t4 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2571 a_8915_n271.t1 a_8902_n286.t3 VSS.t1340 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2572 a_2519_n7203.t0 VCLP.t55 a_2381_n7203.t1 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2573 VSS.t2492 a_4972_4686.t5 a_4877_4671.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2574 VSS.t1428 a_8422_1457.t4 a_8792_1457.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2575 a_7177_437.t1 WWL[13].t16 a_7445_4887.t24 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2576 a_2683_n953.t19 WWLD[4].t13 a_2672_n271.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2577 VSS.t478 a_7272_3425.t4 a_7642_3425.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2578 a_3420_4887.t6 PRE_SRAM.t23 VDD.t2052 VDD.t2051 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2579 a_8902_1201.t0 WWL[10].t15 a_9170_4887.t4 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2580 VSS.t2490 a_372_n271.t5 a_277_n286.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2581 a_4675_n4483.t2 PRE_CLSA.t71 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2582 a_3617_n812.t0 VSS.t635 a_3165_n953.t14 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2583 a_3247_n512.t1 a_3152_n527.t4 VSS.t392 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2584 a_3833_n953.t4 WWL[11].t18 a_3822_975.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2585 VDD.t640 a_6122_693.t5 a_6027_678.t0 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2586 a_4972_975.t1 a_4877_960.t3 VSS.t1703 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2587 a_13171_n8071.t1 Iref3.t13 a_13230_n8026.t1 VSS.t832 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2588 VDD.t511 a_6102_n2234.t3 a_6225_n2132.t1 VDD.t510 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2589 a_2683_n953.t1 WWL[1].t19 a_2672_3425.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2590 a_6708_n953.t5 WWL[12].t16 a_6697_693.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2591 VDD.t13 a_4972_1216.t4 a_4877_1201.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2592 VSS.t1398 a_8993_n2422.t5 a_13602_n4116.t1 VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2593 VSS.t2273 a_372_3425.t5 a_277_3410.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2594 a_742_975.t0 RWLB[11].t10 a_290_n953.t43 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2595 VSS.t328 SAEN.t51 a_11549_n5293.t0 VSS.t304 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2596 a_6697_2421.t1 a_6602_2406.t5 VSS.t1419 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2597 a_1522_1939.t1 a_1427_1924.t3 VDD.t1560 VDD.t1559 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2598 VSS.t2060 a_8997_1216.t3 a_9367_1216.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2599 a_865_n953.t46 RWL[14].t9 a_865_211.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2600 a_8433_n953.t15 WWL[14].t18 a_8422_211.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2601 VSS.t330 SAEN.t52 a_2084_n8026.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2602 a_7858_n953.t2 WWL[8].t15 a_7847_1698.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2603 a_n2642_n6503.t2 a_n2415_n7216.t4 ADC1_OUT[2].t2 VSS.t1416 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2604 a_6040_n512.t0 a_6027_n527.t5 VSS.t1898 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2605 a_6708_n953.t19 WWL[0].t17 a_6697_3666.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2606 a_3042_2662.t1 RWLB[4].t5 a_2590_n953.t36 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2607 a_6697_n271.t1 a_6602_n286.t5 VSS.t231 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2608 a_18_n8071.t0 SAEN.t53 a_215_n8026.t0 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2609 VSS.t490 a_8997_211.t3 a_9367_211.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2610 VDD.t1289 a_4377_n2234.t3 a_4500_n2132.t1 VDD.t1288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2611 a_7858_n953.t12 WWLD[6].t20 a_7847_n812.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2612 a_4315_n953.t44 RWL[4].t6 a_4315_2662.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2613 VDD.t1932 a_8422_975.t4 a_8327_960.t1 VDD.t1931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2614 a_2467_n512.t0 VSS.t634 a_2015_n953.t14 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2615 a_3227_n2234.t0 Din[5].t0 VDD.t860 VDD.t859 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2616 a_2590_n953.t15 VSS.t633 a_2590_4148.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2617 a_8997_4148.t0 a_8902_4133.t4 VSS.t1404 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2618 a_3822_3666.t0 a_3727_3651.t3 VDD.t816 VDD.t815 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2619 VSS.t1574 a_867_n4378.t0 a_867_n4378.t1 VSS.t1573 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2620 a_6697_n30.t1 a_6602_n45.t3 VDD.t1081 VDD.t1080 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2621 a_290_n812.t1 a_277_n827.t5 VSS.t1079 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2622 VDD.t1529 a_372_452.t5 a_277_437.t1 VDD.t1528 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2623 VDD.t634 a_7272_n30.t4 a_7177_n45.t2 VDD.t633 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2624 VDD.t1974 a_7272_n512.t4 a_7177_n527.t2 VDD.t1973 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2625 VDD.t980 a_5857_n5850.t3 ADC8_OUT[1].t1 VDD.t979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2626 VDD.t1890 a_8997_1698.t4 a_8902_1683.t1 VDD.t1889 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2627 VSS.t1608 a_947_n30.t4 a_852_n45.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2628 a_4192_n812.t0 VSS.t632 a_3740_n953.t16 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2629 VDD.t1605 a_7847_3666.t4 a_7752_3651.t0 VDD.t1604 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2630 VSS.t1754 a_947_2662.t5 a_852_2647.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2631 VSS.t1755 a_1522_3184.t4 a_1892_3184.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2632 VDD.t1950 a_372_3666.t4 a_277_3651.t1 VDD.t1949 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2633 a_3493_n4483.t2 ADC6_OUT[0].t3 a_3563_n4470.t2 VSS.t1181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2634 VDD.t1252 a_7252_n2234.t2 a_7375_n2132.t1 VDD.t1251 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2635 SA_OUT[13].t2 a_7785_n1371.t4 a_8028_n1770.t1 VSS.t2034 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2636 a_8422_n812.t2 a_8327_n827.t4 VSS.t1459 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2637 a_2590_3907.t1 a_2577_3892.t5 VSS.t1893 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2638 a_3740_n953.t46 RWL[5].t10 a_3740_2421.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2639 VSS.t2319 a_372_n512.t4 a_742_n512.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2640 VDD.t518 a_8221_n5850.t3 ADC10_OUT[1].t1 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2641 VDD.t1948 a_8997_n812.t4 a_8902_n827.t1 VDD.t1947 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2642 a_4972_3907.t1 a_4877_3892.t4 VDD.t448 VDD.t447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2643 a_6040_n953.t17 RWL[3].t6 a_6040_2943.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2644 a_2097_1457.t1 a_2002_1442.t3 VDD.t600 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2645 VDD.t986 a_7847_693.t5 a_7752_678.t2 VDD.t985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2646 a_n3495_n7203.t0 SAEN.t54 a_n3298_n6847.t0 VSS.t312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2647 a_4890_2943.t1 a_4877_2928.t5 VSS.t930 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2648 a_13934_n4470.t0 SAEN.t55 a_14131_n4114.t0 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2649 a_947_n812.t1 a_852_n827.t4 VSS.t1870 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2650 a_7272_2943.t1 a_7177_2928.t3 VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2651 a_7067_2180.t0 RWLB[6].t7 a_6615_n953.t25 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2652 VDD.t988 a_4397_4686.t4 a_4302_4671.t1 VDD.t987 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2653 a_7283_n953.t21 WWL[0].t18 a_7272_3666.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2654 a_852_2165.t0 WWL[6].t15 a_1120_4887.t22 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2655 a_7858_n953.t5 WWL[10].t16 a_7847_1216.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2656 a_3165_211.t0 a_3152_196.t5 VSS.t939 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2657 a_12963_n7216.t2 ADC14_OUT[2].t3 VDD.t1601 VDD.t1237 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2658 VDD.t1083 a_9405_n8583.t3 ADC11_OUT[3].t1 VDD.t1082 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2659 a_852_437.t2 WWL[13].t17 a_1120_4887.t12 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 a_6615_n953.t44 RWL[13].t7 a_6615_452.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2661 a_5917_n512.t0 VSS.t631 a_5465_n953.t8 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2662 VSS.t1169 a_8422_4686.t4 a_8792_4686.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2663 VSS.t1232 a_2097_2943.t3 a_2467_2943.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2664 VSS.t2083 a_5547_452.t4 a_5452_437.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2665 a_7260_n1770.t1 PRE_VLSA.t26 VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2666 a_8902_4430.t2 WWLD[1].t15 a_9170_4887.t17 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2667 a_3165_3666.t1 a_3152_3651.t5 VSS.t2341 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2668 a_4315_n953.t32 EN.t6 a_4393_n2422.t3 VSS.t1946 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2669 a_4397_452.t1 a_4302_437.t5 VSS.t1315 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2670 a_372_2662.t0 a_277_2647.t4 VSS.t420 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2671 a_9008_n953.t23 WWL[11].t19 a_8997_975.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2672 a_2577_437.t2 WWL[13].t18 a_2845_4887.t22 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2673 a_372_211.t0 a_277_196.t3 VSS.t1033 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2674 a_4890_211.t1 a_4877_196.t5 VSS.t506 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2675 VSS.t2143 a_947_2180.t3 a_1317_2180.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2676 a_7642_n812.t0 VSS.t630 a_7190_n953.t16 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2677 a_7272_n512.t2 a_7177_n527.t4 VSS.t2248 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2678 VDD.t2201 a_4972_4445.t4 a_4877_4430.t2 VDD.t2200 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2679 VDD.t934 a_1522_693.t5 a_1427_678.t2 VDD.t933 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2680 a_2108_n953.t15 WWL[14].t19 a_2097_211.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2681 a_1427_n827.t0 WWLD[6].t21 a_1695_4887.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2682 VSS.t1230 a_8997_4445.t3 a_9367_4445.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2683 a_4315_1939.t1 a_4302_1924.t4 VSS.t819 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2684 VDD.t1809 a_8997_1216.t4 a_8902_1201.t1 VDD.t1808 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2685 a_8422_3907.t1 a_8327_3892.t3 VDD.t1093 VDD.t1092 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2686 a_7765_n953.t33 RWL[7].t11 a_7765_1939.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2687 a_1522_1698.t0 a_1427_1683.t4 VSS.t1442 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2688 VSS.t1073 a_2672_4148.t4 a_2577_4133.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2689 a_5535_n1770.t1 PRE_VLSA.t27 VSS.t124 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2690 VDD.t2054 PRE_SRAM.t24 a_1533_n953.t5 VDD.t2053 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2691 a_6708_n953.t14 WWL[15].t17 a_6697_n30.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2692 a_2590_3425.t1 a_2577_3410.t5 VSS.t235 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2693 a_5547_1939.t1 a_5452_1924.t3 VDD.t806 VDD.t805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2694 a_3833_n953.t18 WWL[14].t20 a_3822_211.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2695 SA_OUT[15].t0 a_8935_n1371.t4 a_9178_n1770.t0 VSS.t978 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2696 a_4972_3425.t2 a_4877_3410.t4 VDD.t940 VDD.t939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2697 a_14072_n8071.t0 VCLP.t56 a_13934_n8071.t1 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2698 VSS.t1770 a_5547_n30.t4 a_5917_n30.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2699 a_3995_4887.t6 PRE_SRAM.t25 a_3833_n953.t5 VDD.t2055 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2700 VSS.t835 a_5547_2943.t3 a_5917_2943.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2701 a_4302_2647.t0 WWL[4].t17 a_4570_4887.t9 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2702 a_7272_693.t2 a_7177_678.t4 VDD.t2142 VDD.t2141 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2703 a_13864_n7216.t1 ADC15_OUT[2].t4 a_13934_n7203.t0 VSS.t1443 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2704 a_5720_4887.t10 WE.t18 a_5768_n2086.t0 VSS.t2391 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2705 a_6615_3666.t1 a_6602_3651.t4 VSS.t1509 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2706 a_8340_n953.t45 RWL[4].t7 a_8340_2662.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2707 a_7765_1698.t1 a_7752_1683.t5 VSS.t2093 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2708 VSS.t1801 a_4397_211.t3 a_4767_211.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2709 a_8221_n7216.t0 PRE_CLSA.t72 VDD.t225 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2710 a_2519_n4470.t0 VCLP.t57 a_2381_n4470.t1 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2711 a_1440_n1053.t1 a_1427_n1068.t5 VSS.t2308 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2712 VSS.t1510 a_4397_1939.t5 a_4302_1924.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2713 a_6492_n512.t1 VSS.t629 a_6040_n953.t16 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2714 a_5917_452.t1 RWLB[13].t10 a_5465_n953.t21 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2715 VDD.t227 PRE_CLSA.t73 ADC10_OUT[1].t0 VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2716 a_865_n953.t44 RWL[4].t8 a_865_2662.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2717 a_2097_1939.t0 a_2002_1924.t5 VSS.t1708 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2718 a_7847_3666.t1 a_7752_3651.t3 VDD.t1593 VDD.t1592 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2719 a_4883_n7203.t0 VCLP.t58 a_4745_n7203.t2 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2720 VSS.t2031 a_4397_2662.t3 a_4767_2662.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2721 VDD.t1806 a_3247_n30.t4 a_3152_n45.t2 VDD.t1805 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2722 a_8410_n1770.t0 PRE_VLSA.t28 VSS.t130 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2723 a_2002_n45.t0 WWL[15].t18 a_2270_4887.t18 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2724 VDD.t229 PRE_CLSA.t74 ADC11_OUT[3].t0 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2725 a_5465_n953.t36 EN.t7 a_5543_n2422.t0 VSS.t1947 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2726 VSS.t1560 a_6697_3184.t5 a_7067_3184.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2727 VDD.t231 PRE_CLSA.t75 ADC8_OUT[3].t0 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2728 a_10797_n5338.t0 VCLP.t59 a_10659_n5338.t1 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2729 a_6122_452.t2 a_6027_437.t3 VSS.t2485 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2730 a_2097_4686.t1 a_2002_4671.t3 VDD.t1564 VDD.t1563 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2731 VSS.t2063 a_4972_2662.t5 a_4877_2647.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2732 a_7247_n7203.t0 a_5743_n6391# a_7109_n7203.t1 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2733 VSS.t2481 a_372_693.t4 a_742_693.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2734 a_n2642_n3770.t2 a_n2415_n4483.t3 ADC1_OUT[0].t1 VSS.t1676 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2735 a_8595_4887.t6 WE.t19 a_8643_n2086.t1 VSS.t2392 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2736 a_7858_n953.t19 WWLD[1].t16 a_7847_4445.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2737 a_4397_3666.t0 a_4302_3651.t5 VSS.t2058 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2738 a_1522_1216.t1 a_1427_1201.t4 VSS.t1531 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2739 a_8422_3425.t1 a_8327_3410.t3 VDD.t1047 VDD.t1046 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2740 VDD.t1352 a_3247_693.t5 a_3152_678.t2 VDD.t1351 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2741 a_1317_1457.t1 RWLB[9].t6 a_865_n953.t28 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2742 VSS.t2324 a_6122_452.t4 a_6492_452.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2743 a_11846_n7203.t1 a_5632_n6430# a_12043_n6847.t0 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2744 VSS.t334 SAEN.t56 a_4448_n8026.t0 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2745 VDD.t398 a_2311_n4483.t4 ADC5_OUT[0].t1 VDD.t397 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2746 VDD.t858 a_2097_2943.t4 a_2002_2928.t1 VDD.t857 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2747 a_6685_n1770.t1 PRE_VLSA.t29 VSS.t128 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2748 a_3727_4133.t2 WWLD[2].t16 a_3995_4887.t17 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2749 a_4877_2165.t2 WWL[6].t16 a_5145_4887.t12 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2750 a_2015_n953.t7 VSS.t628 a_2015_3907.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2751 a_3042_2943.t1 RWLB[3].t5 a_2590_n953.t34 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2752 VDD.t233 PRE_CLSA.t76 ADC1_OUT[3].t0 VDD.t232 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2753 VDD.t235 PRE_CLSA.t77 ADC15_OUT[1].t0 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2754 VSS.t1920 a_6122_2943.t4 a_6492_2943.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2755 a_5547_1939.t0 a_5452_1924.t4 VSS.t1175 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2756 a_7190_3666.t1 a_7177_3651.t5 VSS.t2346 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2757 VDD.t1892 a_947_2180.t4 a_852_2165.t2 VDD.t1891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2758 a_7765_1216.t0 a_7752_1201.t5 VSS.t787 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2759 a_8997_693.t2 a_8902_678.t4 VDD.t740 VDD.t739 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2760 a_6870_4887.t13 WE.t20 a_6918_n2086.t1 VSS.t2393 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 a_3165_n953.t12 VSS.t627 a_3165_n1053.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2762 a_1199_n7203.t0 SAEN.t57 a_1396_n6847.t0 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2763 VSS.t1942 a_4972_2180.t4 a_5342_2180.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2764 VDD.t856 a_8997_4445.t4 a_8902_4430.t0 VDD.t855 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2765 VSS.t1266 a_7847_4148.t5 a_7752_4133.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2766 VSS.t2076 a_8997_2180.t5 a_8902_2165.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2767 VSS.t335 SAEN.t58 a_5630_n5293.t0 VSS.t306 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2768 a_5558_n953.t1 WWL[2].t17 a_5547_3184.t0 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2769 a_8340_1939.t1 a_8327_1924.t5 VSS.t2237 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2770 a_2590_n953.t31 RWL[8].t8 a_2590_1698.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2771 a_8997_1698.t1 a_8902_1683.t4 VSS.t417 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2772 a_n3495_n4470.t0 SAEN.t59 a_n3298_n4114.t0 VSS.t336 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2773 a_1440_n953.t25 RWL[0].t12 a_1440_3666.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2774 a_7847_3666.t0 a_7752_3651.t4 VSS.t1840 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2775 a_13171_n5338.t0 VCLP.t60 a_13033_n5338.t1 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2776 a_865_1939.t0 a_852_1924.t5 VSS.t1646 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2777 a_3727_n45.t0 WWL[15].t19 a_3995_4887.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2778 VDD.t1868 a_10589_n5850.t3 ADC12_OUT[1].t1 VDD.t1508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2779 VDD.t932 a_5547_2943.t4 a_5452_2928.t1 VDD.t931 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2780 VDD.t1392 a_3822_1939.t5 a_3727_1924.t1 VDD.t1391 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2781 a_9170_4887.t23 PRE_SRAM.t26 a_9008_n953.t21 VDD.t2056 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2782 a_3042_693.t1 RWLB[12].t6 a_2590_n953.t20 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2783 a_8327_2165.t2 WWL[6].t17 a_8595_4887.t14 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2784 a_4767_1939.t1 RWLB[7].t11 a_4315_n953.t33 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2785 a_2015_n953.t9 VSS.t626 a_2015_n271.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2786 VSS.t337 SAEN.t60 a_7994_n5293.t0 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2787 a_2590_n953.t9 VSS.t625 a_2590_n812.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2788 a_2672_3184.t1 a_2577_3169.t3 VDD.t1770 VDD.t1769 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2789 a_2672_693.t2 a_2577_678.t4 VDD.t2253 VDD.t2252 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2790 a_7272_n30.t0 a_7177_n45.t3 VSS.t1147 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2791 VSS.t2438 a_n1495_n4378.t6 a_n1495_n4116.t1 VSS.t2433 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2792 VSS.t1968 a_8422_1939.t5 a_8327_1924.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2793 a_3165_n953.t17 RWL[9].t8 a_3165_1457.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2794 a_6122_1457.t0 a_6027_1442.t4 VSS.t1582 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2795 a_2015_n953.t20 RWL[1].t5 a_2015_3425.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2796 VDD.t1786 a_4397_2662.t4 a_4302_2647.t1 VDD.t1785 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2797 a_6615_n953.t7 VSS.t624 a_6615_n1053.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2798 a_4983_n953.t19 WWL[3].t17 a_4972_2943.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2799 VDD.t237 PRE_CLSA.t78 ADC0_OUT[3].t0 VDD.t236 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2800 a_8977_n2234.t0 Din[15].t0 VDD.t1004 VDD.t1003 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2801 VDD.t239 PRE_CLSA.t79 ADC5_OUT[0].t0 VDD.t238 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2802 a_372_2943.t1 a_277_2928.t4 VSS.t768 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2803 VSS.t2075 a_8422_2662.t4 a_8792_2662.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2804 a_8902_2406.t2 WWL[5].t15 a_9170_4887.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2805 a_5465_975.t1 a_5452_960.t5 VSS.t1435 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2806 a_3833_n953.t11 WWL[6].t18 a_3822_2180.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2807 VSS.t2317 a_7843_n2422.t6 a_11514_n4116.t1 VSS.t2312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2808 a_1522_4445.t1 a_1427_4430.t4 VSS.t1127 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2809 a_1522_452.t0 a_1427_437.t4 VSS.t398 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2810 a_8902_n286.t0 WWLD[4].t14 a_9170_4887.t18 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2811 a_902_n6503.t2 VCLP.t61 a_867_n6849.t0 VSS.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2812 VSS.t2180 a_3247_n1053.t5 a_3152_n1068.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2813 a_1317_4686.t0 VSS.t623 a_865_n953.t7 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2814 VDD.t1267 a_4972_2421.t4 a_4877_2406.t2 VDD.t1266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2815 a_8997_1216.t1 a_8902_1201.t4 VSS.t809 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2816 a_2590_n953.t2 RWL[10].t10 a_2590_1216.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2817 VSS.t851 a_8997_2421.t3 a_9367_2421.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2818 a_5342_1457.t0 RWLB[9].t7 a_4890_n953.t36 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2819 VSS.t1660 a_1522_452.t4 a_1892_452.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2820 a_13864_n4483.t1 ADC15_OUT[0].t3 a_13934_n4470.t2 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2821 a_2002_3892.t0 WWLD[3].t19 a_2270_4887.t6 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2822 a_4675_n8583.t2 ADC7_OUT[3].t3 VDD.t1620 VDD.t1619 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2823 VSS.t983 a_6693_n2422.t0 a_6693_n2422.t1 VSS.t982 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2824 a_7765_4445.t1 a_7752_4430.t5 VSS.t1375 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2825 a_4408_n953.t10 WWL[7].t16 a_4397_1939.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2826 a_n52_n8583.t1 ADC3_OUT[3].t3 VDD.t1069 VDD.t1068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2827 a_6040_n953.t8 VSS.t622 a_6040_3907.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2828 a_4302_2928.t0 WWL[3].t18 a_4570_4887.t8 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2829 VSS.t1015 a_2672_1698.t4 a_2577_1683.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2830 a_6615_n953.t18 RWL[9].t9 a_6615_1457.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2831 a_277_4133.t0 WWLD[2].t17 a_545_4887.t17 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2832 a_11549_n5293.t2 a_11776_n5850.t4 ADC13_OUT[1].t2 VSS.t1856 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2833 VDD.t1880 a_7272_4148.t4 a_7177_4133.t1 VDD.t1879 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2834 VDD.t716 a_8422_2180.t4 a_8327_2165.t1 VDD.t715 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2835 VSS.t2194 a_3231_n4378.t6 a_3231_n7825.t1 VSS.t1064 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2836 a_4883_n4470.t0 VCLP.t62 a_4745_n4470.t2 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2837 VDD.t1009 a_3493_n7216.t3 ADC6_OUT[2].t1 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2838 a_4397_693.t2 a_4302_678.t4 VDD.t2116 VDD.t2115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2839 VSS.t339 SAEN.t61 a_n279_n8026.t0 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2840 a_n3357_n5338.t0 VCLP.t63 a_n3495_n5338.t1 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2841 a_7190_n953.t11 VSS.t621 a_7190_n1053.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2842 VSS.t1654 a_2672_n812.t4 a_2577_n827.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2843 VSS.t1241 a_2097_3907.t3 a_2467_3907.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2844 a_n1233_n5850.t2 ADC2_OUT[1].t4 a_n1163_n5338.t2 VSS.t900 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2845 VSS.t1729 a_372_4148.t4 a_742_4148.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2846 VSS.t2074 a_3247_1457.t5 a_3152_1442.t2 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2847 a_9475_n8071.t0 SAEN.t62 a_9672_n8026.t0 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2848 a_7247_n4470.t0 VCLP.t64 a_7109_n4470.t1 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2849 VSS.t1119 a_8997_693.t4 a_8902_678.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2850 a_4890_n953.t10 VSS.t620 a_4890_n512.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 VSS.t1927 a_n314_n4378.t6 a_n314_n7825.t1 VSS.t1924 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2852 VDD.t1457 SA_OUT[4].t3 a_2610_n1371.t1 VDD.t1456 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2853 VDD.t1554 a_n3565_n8583.t3 ADC0_OUT[3].t1 VDD.t1553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2854 a_11846_n4470.t0 SAEN.t63 a_12043_n4114.t0 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2855 a_2519_n4470.t1 Iref0.t5 a_2578_n4114.t1 VSS.t2221 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2856 SA_OUT[11].t2 PRE_VLSA.t30 VDD.t1127 VDD.t1126 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2857 VSS.t2424 a_3822_n1053.t4 a_3727_n1068.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2858 a_2097_n1053.t1 a_2002_n1068.t5 VSS.t896 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2859 VDD.t241 PRE_CLSA.t80 ADC12_OUT[3].t0 VDD.t240 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2860 a_5465_3184.t1 a_5452_3169.t5 VSS.t1653 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2861 a_2097_2662.t1 a_2002_2647.t3 VDD.t341 VDD.t340 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2862 a_5452_3892.t0 WWLD[3].t20 a_5720_4887.t7 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2863 a_8792_1939.t1 RWLB[7].t12 a_8340_n953.t3 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2864 a_6040_n953.t12 VSS.t619 a_6040_n271.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2865 a_3165_n953.t7 VSS.t618 a_3165_4686.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2866 a_6122_4686.t0 a_6027_4671.t4 VSS.t1047 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2867 a_742_3907.t0 VSS.t617 a_290_n953.t17 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2868 VSS.t1445 a_1522_3666.t4 a_1892_3666.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2869 VDD.t850 a_4675_n4483.t4 ADC7_OUT[0].t2 VDD.t849 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2870 a_2577_1924.t0 WWL[7].t17 a_2845_4887.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2871 VSS.t1773 a_1522_n512.t5 a_1427_n527.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2872 a_2002_3410.t0 WWL[1].t20 a_2270_4887.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2873 a_7858_n953.t3 WWL[5].t16 a_7847_2421.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2874 a_2672_n30.t1 a_2577_n45.t4 VSS.t115 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2875 a_1522_n512.t1 a_1427_n527.t4 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2876 a_6040_n953.t21 RWL[1].t6 a_6040_3425.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2877 a_7190_n953.t20 RWL[9].t10 a_7190_1457.t1 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2878 VSS.t1725 a_2672_1216.t4 a_2577_1201.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2879 VSS.t2151 a_2097_n271.t3 a_2467_n271.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2880 a_1199_n4470.t0 SAEN.t64 a_1396_n4114.t0 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2881 a_2015_n812.t1 a_2002_n827.t4 VSS.t1310 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2882 VSS.t1629 a_5547_3907.t3 a_5917_3907.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2883 VDD.t1914 a_2672_n1053.t5 a_2577_n1068.t0 VDD.t1913 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2884 a_3727_1683.t0 WWL[8].t16 a_3995_4887.t21 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2885 VSS.t1627 a_3247_975.t3 a_3617_975.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2886 a_9008_n953.t16 WWL[6].t19 a_8997_2180.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2887 a_865_693.t1 a_852_678.t5 VSS.t2469 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2888 VSS.t820 a_2097_3425.t3 a_2467_3425.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2889 a_3563_n7203.t0 SAEN.t65 a_3760_n6847.t0 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2890 a_3247_n812.t1 a_3152_n827.t3 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2891 a_2590_n953.t7 VSS.t616 a_2590_4445.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2892 a_8997_4445.t1 a_8902_4430.t4 VSS.t2013 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2893 VSS.t876 a_3822_1457.t4 a_3727_1442.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2894 VDD.t502 a_8997_2421.t4 a_8902_2406.t0 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2895 a_9367_693.t0 RWLB[12].t7 a_8915_n953.t42 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2896 a_277_437.t2 WWL[13].t19 a_545_4887.t24 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2897 a_n3565_n4483.t2 ADC0_OUT[0].t4 VDD.t1420 VDD.t1419 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2898 VSS.t1706 a_7272_n1053.t5 a_7177_n1068.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2899 a_5342_4686.t1 VSS.t615 a_4890_n953.t15 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2900 a_5927_n7203.t1 a_5632_n6430# a_6124_n6847.t0 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2901 a_8915_3184.t0 a_8902_3169.t3 VSS.t1237 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2902 a_3740_2180.t0 a_3727_2165.t5 VSS.t990 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2903 a_6122_2180.t2 a_6027_2165.t4 VDD.t1912 VDD.t1911 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2904 a_6615_n953.t2 VSS.t614 a_6615_4686.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2905 VSS.t343 SAEN.t66 a_10362_n5293.t0 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2906 VDD.t1061 SA_OUT[6].t3 a_3760_n1371.t0 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2907 a_3247_n1053.t0 a_3152_n1068.t4 VSS.t2185 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2908 VSS.t1142 a_7847_1698.t5 a_7752_1683.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2909 a_6602_1442.t0 WWL[9].t18 a_6870_4887.t22 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2910 a_5452_3410.t0 WWL[1].t21 a_5720_4887.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2911 a_8433_n953.t14 WWL[7].t18 a_8422_1939.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2912 a_9178_n5293.t2 VCLP.t65 a_9143_n5092.t0 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2913 a_742_3425.t1 RWLB[1].t5 a_290_n953.t27 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2914 a_6615_211.t1 a_6602_196.t4 VSS.t1370 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2915 a_5558_n953.t16 WWL[13].t20 a_5547_452.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2916 VSS.t1107 a_5547_n271.t3 a_5917_n271.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2917 VDD.t870 a_2097_3907.t4 a_2002_3892.t1 VDD.t869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2918 a_958_n953.t8 WWL[7].t19 a_947_1939.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2919 VDD.t371 a_2672_1457.t5 a_2577_1442.t2 VDD.t370 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2920 VSS.t2086 a_7847_n812.t5 a_7752_n827.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2921 a_8221_n5850.t1 ADC10_OUT[1].t3 VDD.t1443 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2922 a_290_n953.t24 RWL[11].t4 a_290_975.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2923 a_n2415_n7216.t1 ADC1_OUT[2].t3 VDD.t1403 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2924 a_1337_n8071.t0 VCLP.t66 a_1199_n8071.t1 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2925 a_n279_n5293.t2 a_n52_n5850.t4 ADC3_OUT[1].t2 VSS.t1251 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2926 VSS.t795 a_3247_4686.t5 a_3152_4671.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2927 VSS.t788 a_6122_3907.t4 a_6492_3907.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2928 a_6697_n812.t1 a_6602_n827.t3 VDD.t1356 VDD.t1355 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2929 VSS.t1017 a_5547_3425.t3 a_5917_3425.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2930 a_7847_452.t1 a_7752_437.t4 VSS.t2448 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2931 a_6697_3184.t1 a_6602_3169.t5 VSS.t1277 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2932 a_3727_1201.t2 WWL[10].t17 a_3995_4887.t8 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2933 VSS.t2376 a_3822_975.t4 a_4192_975.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2934 a_4972_975.t2 a_4877_960.t4 VDD.t1811 VDD.t1810 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2935 a_902_n3770.t1 VCLP.t67 a_867_n4116.t0 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2936 a_5465_n953.t43 RWL[12].t9 a_5465_693.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2937 VSS.t1613 a_7272_1457.t5 a_7177_1442.t0 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2938 VDD.t1360 a_4972_211.t5 a_4877_196.t2 VDD.t1359 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2939 a_11776_n8583.t1 ADC13_OUT[3].t4 a_11846_n8071.t2 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2940 a_6122_n1053.t2 a_6027_n1068.t4 VSS.t1875 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2941 VSS.t2282 a_4397_693.t4 a_4302_678.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2942 a_3266_n6503.t1 VCLP.t68 a_3231_n6849.t0 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2943 a_7190_n953.t48 RWL[14].t10 a_7190_211.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2944 a_6040_n953.t36 EN.t8 a_6268_n2426.t2 VSS.t1948 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2945 VSS.t2348 a_2672_n512.t5 a_3042_n512.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2946 a_3247_n812.t2 a_3152_n827.t4 VSS.t958 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2947 VSS.t1934 a_6697_3666.t5 a_7067_3666.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2948 a_1522_2421.t1 a_1427_2406.t4 VSS.t1349 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2949 a_7752_1924.t2 WWL[7].t20 a_8020_4887.t0 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2950 a_8340_452.t0 a_8327_437.t5 VSS.t923 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2951 VSS.t1261 a_6122_211.t4 a_6027_196.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2952 VDD.t369 a_6697_211.t4 a_6602_196.t0 VDD.t368 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2953 a_n1460_n8026.t2 a_n1233_n8583.t4 ADC2_OUT[3].t2 VSS.t485 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X2954 a_4315_n512.t1 a_4302_n527.t4 VSS.t1603 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2955 a_7190_n953.t9 VSS.t613 a_7190_4686.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2956 a_1317_2662.t1 RWLB[4].t6 a_865_n953.t35 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2957 a_1522_n271.t2 a_1427_n286.t4 VSS.t2089 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2958 VDD.t242 PRE_CLSA.t81 ADC13_OUT[1].t0 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2959 VSS.t945 a_2672_4445.t4 a_2577_4430.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2960 VDD.t1894 a_2097_n271.t4 a_2002_n286.t1 VDD.t1893 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2961 VSS.t793 a_7847_1216.t5 a_7752_1201.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2962 VDD.t1370 a_5547_3907.t4 a_5452_3892.t2 VDD.t1369 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2963 SA_OUT[1].t1 a_885_n1371.t4 a_1128_n1770.t1 VSS.t1930 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2964 a_5547_n512.t1 a_5452_n527.t3 VDD.t1888 VDD.t1887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2965 VDD.t1368 a_3247_975.t4 a_3152_960.t2 VDD.t1367 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2966 a_352_n2234.t0 Din[0].t0 VDD.t872 VDD.t871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2967 VSS.t1027 a_6122_n271.t4 a_6492_n271.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2968 VDD.t488 a_2097_3425.t4 a_2002_3410.t1 VDD.t487 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2969 a_7765_2421.t1 a_7752_2406.t5 VSS.t2059 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2970 a_2683_n953.t14 WWL[15].t20 a_2672_n30.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2971 a_6040_n812.t1 a_6027_n827.t5 VSS.t887 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2972 a_3822_4148.t1 a_3727_4133.t4 VSS.t1072 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2973 a_4972_2180.t1 a_4877_2165.t3 VSS.t1940 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2974 VSS.t1872 a_7272_975.t4 a_7642_975.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2975 VDD.t830 a_6697_n1053.t3 a_6602_n1068.t0 VDD.t829 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2976 a_3740_n953.t1 RWL[2].t12 a_3740_3184.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2977 a_7765_n271.t1 a_7752_n286.t5 VSS.t2291 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2978 VSS.t784 a_5118_n2426.t6 a_5595_n4116.t1 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X2979 VSS.t1389 a_3822_4686.t4 a_3727_4671.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2980 VSS.t1115 a_1522_n30.t3 a_1892_n30.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2981 VSS.t1145 a_6122_3425.t4 a_6492_3425.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2982 a_277_1683.t2 WWL[8].t17 a_545_4887.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2983 a_2270_4887.t24 PRE_SRAM.t27 VDD.t2058 VDD.t2057 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2984 a_4983_n953.t9 WWLD[3].t21 a_4972_3907.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2985 VDD.t777 a_7272_1698.t4 a_7177_1683.t2 VDD.t776 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2986 a_2467_n812.t0 VSS.t612 a_2015_n953.t10 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2987 a_2097_n512.t2 a_2002_n527.t5 VSS.t1995 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2988 a_2683_n953.t23 WWL[11].t20 a_2672_975.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2989 a_5452_n45.t0 WWL[15].t21 a_5720_4887.t20 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2990 VSS.t1353 a_7375_n2132.t2 a_7353_n2086.t1 VSS.t1352 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2991 VSS.t1589 a_372_975.t5 a_277_960.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2992 VSS.t448 a_7847_452.t4 a_8217_452.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2993 a_1129_n7216.t1 ADC4_OUT[2].t3 VDD.t828 VDD.t827 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X2994 a_4767_693.t1 RWLB[12].t8 a_4315_n953.t20 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2995 SA_OUT[6].t1 a_3760_n1371.t4 a_4003_n1770.t1 VSS.t1565 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X2996 a_6602_4671.t0 WWLD[0].t18 a_6870_4887.t7 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2997 VSS.t344 SAEN.t67 a_902_n5293.t0 VSS.t316 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2998 VDD.t1479 a_7272_n812.t4 a_7177_n827.t2 VDD.t1478 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2999 a_4315_n953.t45 RWL[3].t7 a_4315_2943.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3000 a_10659_n8071.t0 SAEN.t68 a_10856_n8026.t0 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3001 a_8997_4148.t1 a_8902_4133.t5 VDD.t1033 VDD.t1032 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3002 VSS.t1846 a_372_1698.t4 a_742_1698.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3003 a_8997_n30.t1 a_8902_n45.t4 VSS.t2255 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3004 a_1533_n953.t14 WWLD[5].t21 a_1522_n512.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3005 a_4883_n4470.t1 Iref0.t6 a_4942_n4114.t1 VSS.t2222 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3006 a_7190_n953.t32 EN.t9 a_7418_n2426.t2 VSS.t1949 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3007 a_6492_211.t0 RWLB[14].t8 a_6040_n953.t41 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3008 VDD.t726 a_5547_n271.t4 a_5452_n286.t1 VDD.t725 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3009 a_4043_n2086.t1 a_3802_n2234.t3 VSS.t847 VSS.t846 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3010 VDD.t1523 a_2672_4686.t5 a_2577_4671.t2 VDD.t1522 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3011 a_5558_n953.t26 WWL[0].t19 a_5547_3666.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3012 a_2097_2943.t2 a_2002_2928.t3 VDD.t1784 VDD.t1783 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3013 a_5630_n5293.t2 a_5857_n5850.t4 ADC8_OUT[1].t2 VSS.t1341 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3014 a_7247_n4470.t1 Iref0.t7 a_7306_n4114.t1 VSS.t2223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3015 VSS.t2018 a_5650_n2132.t2 a_5628_n2086.t1 VSS.t2017 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3016 VSS.t911 a_372_n812.t4 a_742_n812.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3017 VDD.t672 a_5547_3425.t4 a_5452_3410.t2 VDD.t671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3018 a_3165_n953.t26 RWL[4].t9 a_3165_2662.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3019 a_6122_2662.t0 a_6027_2647.t4 VSS.t1557 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3020 VDD.t1632 a_6697_1457.t3 a_6602_1442.t1 VDD.t1631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3021 VDD.t243 PRE_CLSA.t82 ADC7_OUT[2].t0 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3022 a_n1025_n5338.t1 Iref1.t5 a_n966_n5293.t1 VSS.t2224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3023 a_3727_4430.t2 WWLD[1].t17 a_3995_4887.t25 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3024 SA_OUT[3].t1 a_2035_n1371.t4 a_2278_n1770.t0 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3025 VSS.t1373 a_947_2943.t5 a_852_2928.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3026 a_3563_n4470.t0 SAEN.t69 a_3760_n4114.t0 VSS.t346 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3027 VSS.t920 a_7272_4686.t5 a_7177_4671.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3028 a_372_693.t1 a_277_678.t4 VDD.t1994 VDD.t1993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3029 a_4983_n953.t14 WWLD[4].t15 a_4972_n271.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3030 a_7994_n5293.t2 a_8221_n5850.t4 ADC10_OUT[1].t2 VSS.t874 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3031 a_2311_n4483.t2 ADC5_OUT[0].t4 VDD.t1467 VDD.t1466 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3032 VDD.t1125 PRE_VLSA.t31 a_8360_n1371.t2 VDD.t1124 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3033 a_2672_3666.t1 a_2577_3651.t4 VDD.t2094 VDD.t2093 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3034 VSS.t1399 a_8993_n2422.t6 a_13602_n7825.t1 VSS.t1396 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3035 a_5917_n812.t0 VSS.t611 a_5465_n953.t17 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3036 a_5720_4887.t25 PRE_SRAM.t28 VDD.t2060 VDD.t2059 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3037 a_3258_n953.t10 WWL[15].t22 a_3247_n30.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3038 VDD.t1037 a_13864_n7216.t3 ADC15_OUT[2].t1 VDD.t1036 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3039 a_290_n1053.t1 a_277_n1068.t5 VSS.t1192 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3040 a_5547_n512.t2 a_5452_n527.t4 VSS.t2138 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3041 VDD.t1658 a_6122_n512.t4 a_6027_n527.t1 VDD.t1657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3042 a_277_1201.t0 WWL[10].t18 a_545_4887.t5 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3043 a_2015_452.t0 a_2002_437.t4 VSS.t807 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 a_5927_n4470.t0 SAEN.t70 a_6124_n4114.t0 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3045 a_4983_n953.t2 WWL[1].t22 a_4972_3425.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3046 VDD.t1171 a_7272_1216.t4 a_7177_1201.t2 VDD.t1170 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3047 VSS.t1364 a_2097_n30.t4 a_2467_n30.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3048 a_2590_n953.t46 RWL[14].t11 a_2590_211.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3049 VDD.t244 PRE_CLSA.t83 ADC2_OUT[2].t0 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3050 VSS.t1281 a_8525_n2132.t2 a_8503_n2086.t1 VSS.t1280 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3051 a_1510_n1770.t1 PRE_VLSA.t32 VSS.t132 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3052 a_7272_n812.t2 a_7177_n827.t4 VSS.t1719 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3053 VSS.t1308 a_7847_4445.t5 a_7752_4430.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3054 a_2590_n953.t45 RWL[5].t11 a_2590_2421.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3055 a_8997_2421.t1 a_8902_2406.t4 VSS.t1421 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3056 a_3822_1939.t1 a_3727_1924.t4 VDD.t1304 VDD.t1303 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3057 a_947_1457.t1 a_852_1442.t3 VDD.t1827 VDD.t1826 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3058 a_3740_452.t0 a_3727_437.t5 VSS.t1454 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3059 VSS.t1287 a_1522_211.t4 a_1427_196.t0 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3060 a_8997_n271.t1 a_8902_n286.t4 VSS.t2011 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3061 a_8340_n512.t1 a_8327_n527.t5 VSS.t2155 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3062 a_5342_2662.t1 RWLB[4].t7 a_4890_n953.t44 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3063 VSS.t401 a_372_1216.t4 a_742_1216.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3064 a_6122_211.t1 a_6027_196.t4 VDD.t783 VDD.t782 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3065 a_865_n512.t1 a_852_n527.t5 VSS.t1678 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3066 a_13033_n8071.t0 SAEN.t71 a_13230_n8026.t0 VSS.t348 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3067 a_6615_n953.t27 RWL[4].t10 a_6615_2662.t1 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3068 a_1695_4887.t15 WE.t21 a_1743_n2086.t1 VSS.t2394 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3069 a_4767_n512.t0 VSS.t610 a_4315_n953.t13 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3070 a_12736_n8026.t1 VCLP.t69 a_12701_n7825.t0 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3071 VDD.t1656 a_9405_n5850.t3 ADC11_OUT[1].t2 VDD.t1655 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3072 a_4890_n953.t4 VSS.t609 a_4890_4148.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3073 VDD.t1226 a_2097_452.t5 a_2002_437.t1 VDD.t1225 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3074 a_7847_211.t1 a_7752_196.t4 VDD.t974 VDD.t973 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3075 a_3701_n8071.t0 VCLP.t70 a_3563_n8071.t1 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3076 VSS.t2116 a_6800_n2132.t2 a_6778_n2086.t0 VSS.t2115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3077 a_3266_n3770.t1 VCLP.t71 a_3231_n4116.t0 VSS.t177 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3078 a_6492_n1053.t0 VSS.t608 a_6040_n953.t14 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3079 a_6492_n812.t0 VSS.t607 a_6040_n953.t10 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3080 a_8915_975.t0 a_8902_960.t4 VSS.t486 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3081 a_865_n953.t4 RWL[15].t7 a_865_n30.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3082 VSS.t1377 a_3247_2662.t5 a_3152_2647.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3083 VSS.t2099 a_8568_n2426.t5 a_12701_n6849.t1 VSS.t2098 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3084 a_7039_n8583.t0 PRE_CLSA.t84 VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3085 VSS.t1040 a_3247_452.t4 a_3617_452.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3086 a_6065_n8071.t0 VCLP.t72 a_5927_n8071.t1 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3087 a_4890_3907.t1 a_4877_3892.t5 VSS.t771 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3088 a_3165_1939.t0 a_3152_1924.t5 VSS.t1313 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3089 a_2097_975.t1 a_2002_960.t4 VDD.t526 VDD.t525 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3090 a_383_n953.t19 WWLD[7].t17 a_372_n1053.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3091 VSS.t1414 a_1522_4148.t5 a_1427_4133.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3092 a_7272_3907.t1 a_7177_3892.t4 VDD.t1940 VDD.t1939 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3093 VDD.t1210 PRE_A.t8 a_6268_n2426.t3 VDD.t1209 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3094 a_8340_n953.t39 RWL[3].t8 a_8340_2943.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3095 a_4397_1457.t1 a_4302_1442.t3 VDD.t590 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3096 a_9367_2180.t0 RWLB[6].t8 a_8915_n953.t22 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3097 VDD.t866 a_6697_4686.t3 a_6602_4671.t1 VDD.t865 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3098 a_8217_4148.t0 VSS.t606 a_7765_n953.t10 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3099 a_865_n953.t40 RWL[3].t9 a_865_2943.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3100 a_1892_211.t0 RWLB[14].t9 a_1440_n953.t38 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3101 a_977_n1770.t0 a_958_n953.t27 a_935_n1770.t0 VSS.t2178 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3102 a_3152_2165.t2 WWL[6].t20 a_3420_4887.t11 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3103 a_3165_n30.t1 a_3152_n45.t5 VSS.t1971 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3104 a_8997_n1053.t0 a_8902_n1068.t5 VSS.t2270 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3105 a_1317_2943.t0 RWLB[3].t6 a_865_n953.t32 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3106 a_4767_n1053.t0 VSS.t605 a_4315_n953.t4 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3107 VSS.t1356 a_4397_2943.t3 a_4767_2943.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3108 VSS.t1267 a_372_n30.t3 a_742_n30.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3109 a_5465_3666.t0 a_5452_3651.t5 VSS.t2148 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3110 a_7190_n953.t46 RWL[4].t11 a_7190_2662.t1 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3111 VSS.t904 a_2672_2421.t4 a_2577_2406.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3112 VSS.t928 a_4972_2943.t5 a_4877_2928.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3113 a_2845_4887.t26 WE.t22 a_2893_n2086.t0 VSS.t2395 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3114 a_277_4430.t2 WWLD[1].t18 a_545_4887.t18 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3115 VSS.t387 a_3247_2180.t3 a_3617_2180.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3116 a_372_n30.t0 a_277_n45.t4 VSS.t981 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3117 a_4890_n30.t0 a_4877_n45.t5 VSS.t1490 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3118 VDD.t385 a_7272_4445.t4 a_7177_4430.t2 VDD.t384 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3119 a_5857_n8583.t2 ADC8_OUT[3].t4 a_5927_n8071.t2 VSS.t800 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3120 VDD.t1212 PRE_A.t9 a_8993_n2422.t3 VDD.t1211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3121 a_7752_678.t0 WWL[12].t17 a_8020_4887.t14 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3122 VSS.t1158 a_6268_n2426.t6 a_7959_n4116.t1 VSS.t1153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3123 a_383_n953.t20 WWL[9].t19 a_372_1457.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 VSS.t1068 a_3822_2662.t4 a_3727_2647.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3125 a_6615_1939.t1 a_6602_1924.t4 VSS.t1381 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3126 a_3822_1698.t2 a_3727_1683.t4 VSS.t2147 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3127 a_9405_n7216.t0 PRE_CLSA.t85 VDD.t247 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3128 VSS.t2134 a_7418_n2426.t6 a_10327_n4116.t1 VSS.t2129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3129 a_7642_n1053.t0 VSS.t604 a_7190_n953.t10 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3130 a_947_4686.t2 a_852_4671.t3 VDD.t810 VDD.t809 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3131 VDD.t2062 PRE_SRAM.t29 a_3833_n953.t6 VDD.t2061 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3132 a_n2642_n6503.t1 VCLP.t73 a_n2677_n6849.t0 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3133 VDD.t248 PRE_CLSA.t86 ADC11_OUT[1].t0 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3134 VSS.t2337 a_372_4445.t4 a_742_4445.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3135 a_7847_1939.t1 a_7752_1924.t3 VDD.t1644 VDD.t1643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3136 VDD.t249 PRE_CLSA.t87 ADC8_OUT[1].t0 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3137 a_4890_3425.t1 a_4877_3410.t5 VSS.t1304 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3138 a_7272_3425.t1 a_7177_3410.t4 VDD.t1388 VDD.t1387 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3139 a_13637_n6503.t2 a_5743_n6391# a_13602_n6849.t0 VSS.t200 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3140 a_4960_n1770.t1 a_5145_4887.t27 a_5153_n1770.t0 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3141 VDD.t1214 PRE_A.t10 a_7418_n2426.t3 VDD.t1213 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3142 a_6602_2647.t0 WWL[4].t18 a_6870_4887.t23 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3143 a_1522_211.t1 a_1427_196.t4 VDD.t1666 VDD.t1665 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3144 a_8902_3169.t0 WWL[2].t18 a_9170_4887.t24 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3145 a_7067_975.t0 RWLB[11].t11 a_6615_n953.t24 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3146 a_8915_3666.t0 a_8902_3651.t3 VSS.t1216 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3147 VSS.t1808 a_6697_1939.t4 a_6602_1924.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3148 a_8792_n512.t0 VSS.t603 a_8340_n953.t10 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3149 VDD.t568 a_2672_2662.t5 a_2577_2647.t1 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3150 a_8997_1698.t2 a_8902_1683.t5 VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3151 a_4397_1939.t1 a_4302_1924.t5 VSS.t1188 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3152 SA_OUT[12].t1 a_7210_n1371.t3 VDD.t1798 VDD.t1797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3153 a_5917_n1053.t0 VSS.t602 a_5465_n953.t13 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3154 a_2577_n527.t0 WWLD[5].t22 a_2845_4887.t5 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3155 VDD.t377 a_4972_3184.t4 a_4877_3169.t2 VDD.t376 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3156 a_6122_2943.t1 a_6027_2928.t4 VSS.t817 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3157 a_290_n953.t32 RWL[6].t5 a_290_2180.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3158 a_10362_n5293.t2 a_10589_n5850.t4 ADC12_OUT[1].t2 VSS.t1815 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3159 VDD.t250 PRE_CLSA.t88 ADC1_OUT[1].t0 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3160 a_8792_975.t0 RWLB[11].t12 a_8340_n953.t40 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3161 VSS.t1074 a_2672_4148.t5 a_3042_4148.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3162 VSS.t1205 a_8997_3184.t3 a_9367_3184.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3163 VSS.t425 a_3822_2180.t4 a_4192_2180.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3164 a_6812_n6503.t0 a_7039_n7216.t4 ADC9_OUT[2].t2 VSS.t991 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3165 a_3727_2406.t2 WWL[5].t17 a_3995_4887.t12 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3166 a_7835_n1770.t1 a_8020_4887.t27 a_8028_n1770.t0 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3167 a_4397_4686.t1 a_4302_4671.t3 VDD.t1607 VDD.t1606 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3168 VSS.t419 a_7272_2662.t5 a_7177_2647.t0 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3169 a_3727_n286.t0 WWLD[4].t16 a_3995_4887.t16 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3170 a_6697_3666.t0 a_6602_3651.t5 VSS.t1180 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3171 a_7190_1939.t1 a_7177_1924.t5 VSS.t1701 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3172 a_7039_n4483.t2 ADC9_OUT[0].t4 VDD.t1254 VDD.t1253 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3173 a_3822_1216.t2 a_3727_1201.t4 VSS.t1722 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3174 SA_OUT[9].t0 a_5485_n1371.t3 VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3175 a_3247_452.t2 a_3152_437.t4 VDD.t1804 VDD.t1803 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3176 a_3042_3907.t0 VSS.t601 a_2590_n953.t8 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3177 VDD.t992 a_4397_2943.t4 a_4302_2928.t1 VDD.t991 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3178 a_3617_1457.t1 RWLB[9].t8 a_3165_n953.t33 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3179 a_7177_2165.t0 WWL[6].t21 a_7445_4887.t13 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3180 a_6027_4133.t0 WWLD[2].t18 a_6295_4887.t14 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3181 a_5342_2943.t1 RWLB[3].t7 a_4890_n953.t41 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3182 a_4315_n953.t12 VSS.t600 a_4315_3907.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3183 VSS.t2126 a_8422_2943.t4 a_8792_2943.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3184 VSS.t891 a_7847_2421.t5 a_7752_2406.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3185 a_6110_n1770.t0 a_6295_4887.t27 a_6303_n1770.t0 VSS.t1511 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3186 a_2015_n953.t21 RWL[11].t5 a_2015_975.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3187 VDD.t1583 a_8422_452.t5 a_8327_437.t2 VDD.t1582 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3188 VDD.t319 a_3247_2180.t4 a_3152_2165.t0 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3189 a_7847_1939.t0 a_7752_1924.t4 VSS.t1881 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3190 a_8997_1216.t2 a_8902_1201.t5 VDD.t478 VDD.t477 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3191 a_5465_n953.t5 VSS.t599 a_5465_n1053.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3192 VSS.t2474 a_7272_2180.t4 a_7642_2180.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3193 a_n2207_n8071.t1 Iref3.t14 a_n2148_n8026.t1 VSS.t1978 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3194 a_383_n953.t6 WWLD[0].t19 a_372_4686.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3195 VSS.t349 SAEN.t72 a_9178_n5293.t0 VSS.t323 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3196 SA_OUT[14].t1 a_8360_n1371.t3 VDD.t1236 VDD.t1235 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3197 VSS.t870 a_947_3907.t5 a_852_3892.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3198 a_8422_975.t1 a_8327_960.t4 VDD.t1924 VDD.t1923 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3199 a_3152_678.t0 WWL[12].t18 a_3420_4887.t10 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3200 VSS.t351 SAEN.t73 a_n1460_n8026.t0 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3201 a_8915_n953.t31 RWL[12].t10 a_8915_693.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3202 VDD.t251 PRE_CLSA.t89 ADC0_OUT[1].t0 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3203 VDD.t2064 PRE_SRAM.t30 a_9008_n953.t22 VDD.t2063 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3204 a_1533_n953.t17 WWLD[2].t19 a_1522_4148.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3205 a_7858_n953.t26 WWL[2].t19 a_7847_3184.t0 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3206 a_2683_n953.t16 WWL[6].t22 a_2672_2180.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3207 VSS.t1334 a_7847_211.t4 a_7752_196.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3208 a_3740_n953.t0 RWL[0].t13 a_3740_3666.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3209 VSS.t471 a_372_2180.t5 a_277_2165.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3210 a_4890_n953.t37 RWL[8].t9 a_4890_1698.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 VSS.t352 SAEN.t74 a_2084_n6503.t0 VSS.t329 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3212 a_4877_196.t0 WWL[14].t21 a_5145_4887.t17 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3213 a_8985_n1770.t2 a_9170_4887.t27 a_9178_n1770.t1 VSS.t2187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3214 VSS.t1379 a_2097_n1053.t5 a_2002_n1068.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3215 a_6697_693.t1 a_6602_678.t5 VSS.t1100 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3216 VSS.t2439 a_n1495_n4378.t7 a_n1495_n7825.t1 VSS.t2436 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3217 SA_OUT[4].t2 PRE_VLSA.t33 VDD.t1123 VDD.t1122 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3218 VSS.t1218 a_7847_1939.t3 a_8217_1939.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3219 a_290_1457.t1 a_277_1442.t5 VSS.t915 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3220 a_18_n7203.t0 SAEN.t75 a_215_n6847.t0 VSS.t331 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3221 a_4315_n953.t16 VSS.t598 a_4315_n271.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3222 a_4890_n953.t3 VSS.t597 a_4890_n812.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3223 a_4192_1457.t1 RWLB[9].t9 a_3740_n953.t30 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3224 SA_OUT[11].t0 a_6635_n1371.t3 VDD.t572 VDD.t571 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3225 a_545_4887.t23 PRE_SRAM.t31 a_383_n953.t4 VDD.t2065 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3226 a_3042_3425.t0 RWLB[1].t6 a_2590_n953.t27 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3227 a_n1163_n5338.t0 SAEN.t76 a_n966_n5293.t0 VSS.t325 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3228 a_3258_n953.t6 WWL[7].t21 a_3247_1939.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3229 VSS.t1826 a_1522_1698.t5 a_1427_1683.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3230 a_2467_975.t0 RWLB[11].t13 a_2015_n953.t41 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3231 a_7752_n527.t0 WWLD[5].t23 a_8020_4887.t3 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3232 a_4315_n953.t21 RWL[1].t7 a_4315_3425.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3233 a_5465_n953.t19 RWL[9].t11 a_5465_1457.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3234 a_8422_1457.t0 a_8327_1442.t4 VSS.t1113 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3235 a_8915_n953.t4 VSS.t596 a_8915_n1053.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3236 VDD.t2120 a_6697_2662.t3 a_6602_2647.t1 VDD.t2119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 VSS.t353 SAEN.t77 a_n2642_n5293.t0 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3238 VDD.t2227 a_6122_4148.t4 a_6027_4133.t2 VDD.t2226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3239 a_372_3907.t2 a_277_3892.t4 VSS.t2260 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3240 VDD.t836 a_8997_3184.t4 a_8902_3169.t1 VDD.t835 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3241 a_8217_1698.t1 RWLB[8].t10 a_7765_n953.t35 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3242 a_947_1457.t0 a_852_1442.t4 VSS.t2079 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3243 a_7190_693.t1 a_7177_678.t5 VSS.t2344 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3244 VSS.t2318 a_7843_n2422.t7 a_11514_n7825.t1 VSS.t2315 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3245 a_4675_n5850.t1 ADC7_OUT[1].t3 VDD.t1571 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3246 a_n52_n5850.t1 ADC3_OUT[1].t3 VDD.t743 VDD.t681 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3247 VSS.t1568 a_947_n271.t5 a_852_n286.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3248 VSS.t1463 a_1522_n812.t5 a_1427_n827.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3249 a_1522_n812.t2 a_1427_n827.t4 VDD.t524 VDD.t523 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3250 a_3822_4445.t1 a_3727_4430.t4 VSS.t1054 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3251 VSS.t1680 a_2097_1457.t5 a_2002_1442.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3252 a_n2642_n3770.t1 VCLP.t74 a_n2677_n4116.t0 VSS.t180 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3253 VSS.t1804 a_947_3425.t5 a_852_3410.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3254 a_277_2406.t0 WWL[5].t18 a_545_4887.t3 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3255 a_8217_211.t1 RWLB[14].t10 a_7765_n953.t47 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3256 a_n1025_n7203.t1 Iref2.t5 a_n966_n6847.t1 VSS.t1983 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3257 VSS.t1997 a_5547_n1053.t5 a_5452_n1068.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3258 a_3617_4686.t0 VSS.t595 a_3165_n953.t2 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3259 VDD.t2180 a_7272_2421.t4 a_7177_2406.t1 VDD.t2179 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3260 a_947_452.t2 a_852_437.t5 VSS.t2432 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3261 a_277_n286.t2 WWLD[4].t17 a_545_4887.t9 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3262 a_10589_n8583.t2 ADC12_OUT[3].t4 a_10659_n8071.t2 VSS.t1530 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3263 a_13637_n3770.t1 VCLP.t75 a_13602_n4116.t0 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3264 a_4890_n953.t35 RWL[10].t11 a_4890_1216.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3265 a_6133_n953.t15 WWL[12].t19 a_6122_693.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3266 a_7642_1457.t1 RWLB[9].t10 a_7190_n953.t28 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3267 a_4302_3892.t0 WWLD[3].t22 a_4570_4887.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3268 a_947_2662.t1 a_852_2647.t3 VDD.t755 VDD.t754 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3269 a_6708_n953.t8 WWL[7].t22 a_6697_1939.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3270 a_1427_1442.t2 WWL[9].t20 a_1695_4887.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3271 a_8340_n953.t15 VSS.t594 a_8340_3907.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3272 VSS.t1674 a_372_2421.t4 a_742_2421.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3273 a_8915_n953.t35 RWL[9].t12 a_8915_1457.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3274 VSS.t1087 a_6697_693.t5 a_7067_693.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3275 a_8422_693.t0 a_8327_678.t4 VSS.t894 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3276 a_290_n953.t1 RWL[14].t12 a_290_211.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3277 VDD.t363 a_n3565_n5850.t3 ADC0_OUT[1].t2 VDD.t362 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3278 a_8997_4445.t2 a_8902_4430.t5 VDD.t1067 VDD.t1066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3279 a_6602_2928.t2 WWL[3].t19 a_6870_4887.t20 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3280 a_6040_n953.t24 RWL[11].t6 a_6040_975.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3281 VDD.t252 PRE_CLSA.t90 ADC12_OUT[1].t0 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3282 VDD.t1101 a_3822_452.t4 a_3727_437.t1 VDD.t1100 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3283 a_865_n953.t10 VSS.t593 a_865_3907.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3284 VSS.t1553 a_1522_1216.t5 a_1427_1201.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3285 a_12963_n7216.t1 ADC14_OUT[2].t4 a_13033_n7203.t2 VSS.t1540 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3286 a_6812_n3770.t1 a_7039_n4483.t3 ADC9_OUT[0].t1 VSS.t429 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3287 VSS.t1469 a_4397_3907.t3 a_4767_3907.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3288 a_372_3425.t2 a_277_3410.t4 VSS.t2276 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3289 a_8217_1216.t1 RWLB[10].t10 a_7765_n953.t45 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3290 VSS.t1412 a_8422_693.t4 a_8792_693.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3291 VDD.t1952 a_1522_n1053.t4 a_1427_n1068.t0 VDD.t1951 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3292 a_1522_3184.t0 a_1427_3169.t4 VSS.t1566 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3293 VSS.t1780 a_2097_975.t3 a_2467_975.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3294 a_4315_n953.t1 RWL[14].t13 a_4315_211.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3295 VSS.t1749 a_4972_3907.t5 a_4877_3892.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3296 VSS.t1687 a_5547_1457.t5 a_5452_1442.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3297 a_3822_975.t1 a_3727_960.t4 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3298 a_14072_n5338.t1 Iref1.t6 a_14131_n5293.t1 VSS.t2225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3299 a_290_4686.t1 a_277_4671.t5 VSS.t1528 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3300 VDD.t842 a_7847_1939.t4 a_7752_1924.t0 VDD.t841 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3301 VSS.t1598 a_3247_211.t4 a_3152_196.t2 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3302 a_n279_n5293.t1 VCLP.t76 a_n314_n5092.t0 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3303 a_2097_211.t0 a_2002_196.t5 VSS.t1258 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3304 VSS.t1225 a_947_n512.t3 a_1317_n512.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3305 a_4192_4686.t0 VSS.t592 a_3740_n953.t6 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3306 VSS.t1864 a_6122_n1053.t5 a_6027_n1068.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3307 VDD.t404 a_372_1939.t4 a_277_1924.t1 VDD.t403 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3308 VSS.t1016 a_2672_1698.t5 a_3042_1698.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3309 a_8221_n5850.t2 ADC10_OUT[1].t4 a_8291_n5338.t2 VSS.t1698 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3310 a_1440_4148.t1 a_1427_4133.t5 VSS.t1845 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3311 a_7765_3184.t0 a_7752_3169.t5 VSS.t806 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3312 a_4397_2662.t1 a_4302_2647.t3 VDD.t854 VDD.t853 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3313 a_2590_2180.t0 a_2577_2165.t5 VSS.t1525 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3314 a_4972_2180.t2 a_4877_2165.t4 VDD.t1714 VDD.t1713 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3315 a_7190_n953.t3 RWL[15].t8 a_7190_n30.t1 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3316 a_8340_n953.t9 VSS.t591 a_8340_n271.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3317 a_5465_n953.t7 VSS.t590 a_5465_4686.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3318 a_8422_4686.t1 a_8327_4671.t4 VSS.t1401 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3319 a_865_n953.t9 VSS.t589 a_865_n271.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3320 VSS.t2457 a_2049_n4378.t5 a_2049_n6849.t1 VSS.t2456 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3321 VSS.t1655 a_2672_n812.t5 a_3042_n812.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3322 a_947_4686.t1 a_852_4671.t4 VSS.t1178 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3323 a_4302_3410.t0 WWL[1].t23 a_4570_4887.t3 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3324 a_7283_n953.t9 WWL[7].t23 a_7272_1939.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3325 a_3822_n512.t2 a_3727_n527.t4 VDD.t2182 VDD.t2181 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3326 a_8340_n953.t25 RWL[1].t8 a_8340_3425.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3327 VSS.t1880 a_4397_n271.t3 a_4767_n271.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3328 a_12963_n7216.t0 PRE_CLSA.t91 VDD.t253 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3329 VDD.t834 a_1522_1457.t4 a_1427_1442.t1 VDD.t833 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3330 a_6040_n953.t42 RWL[13].t8 a_6040_452.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3331 a_4315_n812.t1 a_4302_n827.t4 VSS.t2239 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3332 a_865_n953.t24 RWL[1].t9 a_865_3425.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3333 VSS.t772 a_5547_975.t3 a_5917_975.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3334 a_2590_693.t1 a_2577_678.t5 VSS.t2499 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3335 a_6027_1683.t2 WWL[8].t18 a_6295_4887.t22 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3336 VSS.t1824 a_4972_n271.t5 a_4877_n286.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3337 VSS.t840 a_2097_4686.t5 a_2002_4671.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3338 VSS.t1544 a_4972_452.t4 a_4877_437.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3339 VDD.t1831 a_5547_452.t5 a_5452_437.t1 VDD.t1830 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3340 a_5547_n812.t1 a_5452_n827.t3 VDD.t1722 VDD.t1721 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3341 VSS.t2029 a_4397_3425.t3 a_4767_3425.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3342 VSS.t355 SAEN.t78 a_2084_n3770.t0 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3343 a_4890_n953.t2 VSS.t588 a_4890_4445.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3344 a_2108_n953.t19 WWLD[7].t18 a_2097_n1053.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3345 VSS.t1306 a_4972_3425.t5 a_4877_3410.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3346 a_383_n953.t21 WWL[4].t19 a_372_2662.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3347 VSS.t966 a_6122_1457.t5 a_6027_1442.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3348 a_7642_4686.t0 VSS.t587 a_7190_n953.t12 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3349 a_3617_211.t0 RWLB[14].t11 a_3165_n953.t41 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3350 VDD.t556 a_352_n2234.t3 a_475_n2132.t1 VDD.t555 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3351 VSS.t356 SAEN.t79 a_4448_n6503.t0 VSS.t333 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3352 a_11549_n6503.t1 a_5743_n6391# a_11514_n6849.t1 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3353 a_18_n4470.t0 SAEN.t80 a_215_n4114.t0 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3354 VDD.t1121 PRE_VLSA.t34 a_1460_n1371.t0 VDD.t1120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3355 a_1427_4671.t0 WWLD[0].t20 a_1695_4887.t7 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3356 a_8422_2180.t1 a_8327_2165.t4 VDD.t718 VDD.t717 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3357 a_8915_n953.t7 VSS.t586 a_8915_4686.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3358 a_1533_n953.t10 WWL[12].t20 a_1522_693.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3359 a_6102_n2234.t1 Din[10].t1 VSS.t1369 VSS.t1368 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3360 a_2097_n812.t2 a_2002_n827.t5 VSS.t1441 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3361 VSS.t1726 a_2672_1216.t5 a_3042_1216.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3362 a_1533_n953.t21 WWL[8].t19 a_1522_1698.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3363 a_3165_n512.t1 a_3152_n527.t5 VSS.t400 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3364 VSS.t1523 a_1522_4445.t5 a_1427_4430.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3365 VSS.t943 a_2097_693.t4 a_2467_693.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3366 a_6615_n30.t0 a_6602_n45.t4 VSS.t1438 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3367 a_902_n8026.t2 a_1129_n8583.t4 ADC4_OUT[3].t2 VSS.t1045 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3368 a_3822_693.t0 a_3727_678.t5 VSS.t250 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3369 a_360_n1770.t1 PRE_VLSA.t35 VSS.t134 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3370 a_8217_4445.t0 VSS.t585 a_7765_n953.t8 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3371 VDD.t1189 a_4397_3907.t4 a_4302_3892.t1 VDD.t1188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3372 VSS.t1999 a_1625_n2132.t2 a_1603_n2086.t0 VSS.t1998 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3373 a_1533_n953.t1 WWLD[6].t22 a_1522_n812.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3374 VDD.t1527 a_2097_975.t4 a_2002_960.t2 VDD.t1526 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3375 a_7177_960.t0 WWL[11].t21 a_7445_4887.t23 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3376 SA_OUT[9].t2 PRE_VLSA.t36 VDD.t1119 VDD.t1118 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3377 VSS.t415 a_5547_4686.t5 a_5452_4671.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3378 VSS.t412 a_8422_3907.t4 a_8792_3907.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3379 VSS.t1507 a_3822_211.t4 a_4192_211.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3380 VDD.t1117 PRE_VLSA.t37 a_4335_n1371.t2 VDD.t1116 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3381 a_2672_4148.t2 a_2577_4133.t4 VSS.t1515 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3382 a_2590_n953.t1 RWL[2].t13 a_2590_3184.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3383 a_8997_3184.t1 a_8902_3169.t4 VSS.t1238 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3384 VSS.t2470 a_6122_975.t4 a_6492_975.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3385 a_8902_3651.t2 WWL[0].t20 a_9170_4887.t16 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3386 a_2108_n953.t20 WWL[9].t21 a_2097_1457.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3387 a_6027_1201.t0 WWL[10].t19 a_6295_4887.t7 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3388 a_5342_452.t1 RWLB[13].t11 a_4890_n953.t20 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3389 VSS.t1006 a_7272_n30.t5 a_7177_n45.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3390 VDD.t976 a_947_n512.t4 a_852_n527.t1 VDD.t975 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3391 VDD.t391 a_4972_3666.t4 a_4877_3651.t1 VDD.t390 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3392 VDD.t530 a_6122_1698.t4 a_6027_1683.t1 VDD.t529 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3393 a_n1025_n8071.t0 VCLP.t77 a_n1163_n8071.t1 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3394 VSS.t1109 a_4972_n512.t4 a_5342_n512.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 a_156_n8071.t0 VCLP.t78 a_18_n8071.t1 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3396 a_5547_n812.t2 a_5452_n827.t4 VSS.t1960 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3397 VSS.t1625 a_8997_3666.t3 a_9367_3666.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3398 a_3822_2421.t1 a_3727_2406.t4 VSS.t913 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3399 SA_OUT[14].t0 PRE_VLSA.t38 VDD.t1115 VDD.t1114 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3400 VDD.t1326 a_6122_n812.t4 a_6027_n827.t2 VDD.t1325 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3401 a_3165_n953.t16 RWL[3].t10 a_3165_2943.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3402 VSS.t1741 a_8997_n512.t5 a_8902_n527.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3403 a_6615_n512.t1 a_6602_n527.t4 VSS.t2509 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3404 a_3617_2662.t0 RWLB[4].t8 a_3165_n953.t39 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3405 a_3822_n271.t1 a_3727_n286.t4 VSS.t1383 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3406 VDD.t1113 PRE_VLSA.t39 a_2610_n1371.t0 VDD.t1112 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3407 a_947_2943.t2 a_852_2928.t3 VDD.t922 VDD.t921 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3408 VDD.t1314 a_4397_n271.t4 a_4302_n286.t2 VDD.t1313 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3409 a_7252_n2234.t0 Din[12].t1 VSS.t1691 VSS.t1690 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3410 VDD.t1380 a_1522_4686.t4 a_1427_4671.t2 VDD.t1379 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3411 a_372_4148.t0 a_277_4133.t4 VDD.t958 VDD.t957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3412 a_7847_n512.t1 a_7752_n527.t3 VDD.t1487 VDD.t1486 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3413 a_1533_n953.t8 WWL[10].t20 a_1522_1216.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3414 VDD.t460 a_5547_975.t4 a_5452_960.t1 VDD.t459 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3415 VSS.t785 a_5118_n2426.t7 a_5595_n7825.t1 VSS.t782 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3416 a_12963_n4483.t1 ADC14_OUT[0].t3 a_13033_n4470.t2 VSS.t1484 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3417 VDD.t1216 PRE_A.t11 a_n2677_n4378.t3 VDD.t1215 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3418 a_1892_4148.t0 VSS.t584 a_1440_n953.t10 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3419 a_2015_n953.t30 RWL[6].t6 a_2015_2180.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3420 VSS.t2009 a_8422_n271.t4 a_8792_n271.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3421 a_8340_n812.t1 a_8327_n827.t5 VSS.t1460 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3422 VDD.t1260 a_4397_3425.t4 a_4302_3410.t1 VDD.t1259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3423 a_8997_2421.t2 a_8902_2406.t5 VDD.t1051 VDD.t1050 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3424 a_1440_n953.t39 RWL[13].t9 a_1440_452.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3425 a_n3357_n5338.t1 Iref1.t7 a_n3298_n5293.t1 VSS.t2226 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3426 a_2672_n1053.t1 a_2577_n1068.t5 VDD.t2144 VDD.t2143 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3427 a_865_n812.t1 a_852_n827.t5 VSS.t1871 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3428 VSS.t1279 a_6122_4686.t5 a_6027_4671.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3429 VSS.t1004 a_8422_3425.t4 a_8792_3425.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3430 a_8997_n271.t2 a_8902_n286.t5 VDD.t1774 VDD.t1773 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3431 a_4570_4887.t21 PRE_SRAM.t32 VDD.t2067 VDD.t2066 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3432 a_4767_n812.t0 VSS.t583 a_4315_n953.t15 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3433 a_4397_n512.t2 a_4302_n527.t5 VSS.t1604 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3434 a_4983_n953.t4 WWL[11].t22 a_4972_975.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3435 a_6602_196.t1 WWL[14].t22 a_6870_4887.t17 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3436 VDD.t1111 PRE_VLSA.t40 a_5485_n1371.t0 VDD.t1110 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3437 a_6133_n953.t26 WWLD[7].t19 a_6122_n1053.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3438 VSS.t1645 a_7847_n30.t5 a_7752_n45.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3439 VSS.t946 a_2672_4445.t5 a_3042_4445.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3440 VDD.t796 a_6122_1216.t4 a_6027_1201.t1 VDD.t795 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3441 a_2097_3907.t1 a_2002_3892.t3 VDD.t1874 VDD.t1873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3442 VSS.t2021 a_2672_3184.t4 a_2577_3169.t1 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3443 a_6615_n953.t17 RWL[3].t11 a_6615_2943.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3444 a_1440_n953.t27 RWL[7].t12 a_1440_1939.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3445 a_9178_n5293.t1 a_9405_n5850.t4 ADC11_OUT[1].t1 VSS.t1386 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3446 VDD.t1218 PRE_A.t12 a_n314_n4378.t3 VDD.t1217 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3447 a_8503_n2086.t0 WE.t23 a_8433_n953.t12 VSS.t2396 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3448 a_290_2662.t0 a_277_2647.t5 VSS.t421 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3449 a_3833_n953.t13 WWLD[5].t24 a_3822_n512.t1 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3450 a_4397_2943.t2 a_4302_2928.t3 VDD.t868 VDD.t867 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3451 a_2672_1939.t2 a_2577_1924.t4 VDD.t1589 VDD.t1588 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3452 a_852_960.t0 WWL[11].t23 a_1120_4887.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3453 a_6697_452.t0 a_6602_437.t4 VDD.t1017 VDD.t1016 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3454 a_6492_n30.t1 RWLB[15].t9 a_6040_n953.t37 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3455 a_7858_n953.t21 WWL[0].t21 a_7847_3666.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3456 a_4972_n1053.t0 a_4877_n1068.t4 VSS.t2366 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3457 a_7190_n512.t1 a_7177_n527.t5 VSS.t2236 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3458 a_4192_2662.t0 RWLB[4].t9 a_3740_n953.t36 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3459 a_5547_n1053.t1 a_5452_n1068.t5 VDD.t444 VDD.t443 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3460 VSS.t358 SAEN.t81 a_n279_n6503.t0 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3461 a_5465_n953.t47 RWL[4].t12 a_5465_2662.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3462 a_8422_2662.t0 a_8327_2647.t4 VSS.t1918 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3463 a_1440_1698.t1 a_1427_1683.t5 VSS.t1309 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3464 a_4397_975.t2 a_4302_960.t5 VSS.t2108 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3465 a_2108_n953.t8 WWLD[0].t21 a_2097_4686.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3466 a_6027_4430.t2 WWLD[1].t19 a_6295_4887.t23 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3467 VSS.t1003 a_3247_2943.t5 a_3152_2928.t2 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3468 a_947_2662.t0 a_852_2647.t4 VSS.t867 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3469 a_2577_960.t0 WWL[11].t24 a_2845_4887.t21 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3470 a_9475_n7203.t1 a_5632_n6430# a_9672_n6847.t0 VSS.t340 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3471 a_7847_n512.t2 a_7752_n527.t4 VSS.t1742 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3472 a_6133_n953.t14 WWL[9].t22 a_6122_1457.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3473 VDD.t614 a_8422_n512.t4 a_8327_n527.t1 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3474 a_3266_n6503.t2 a_3493_n7216.t4 ADC6_OUT[2].t2 VSS.t1376 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3475 a_7858_n953.t7 WWL[12].t21 a_7847_693.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3476 a_11549_n3770.t2 VCLP.t79 a_11514_n4116.t0 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3477 VSS.t360 SAEN.t82 a_4448_n3770.t0 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3478 a_3822_n1053.t2 a_3727_n1068.t5 VDD.t2215 VDD.t2214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3479 VDD.t1366 a_8997_3666.t4 a_8902_3651.t0 VDD.t1365 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3480 VSS.t1513 a_2097_2662.t5 a_2002_2647.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3481 VDD.t255 PRE_CLSA.t92 ADC14_OUT[3].t0 VDD.t254 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3482 a_2015_1457.t0 a_2002_1442.t4 VSS.t954 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3483 a_4890_n953.t34 RWL[5].t12 a_4890_2421.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3484 a_3493_n4483.t1 ADC6_OUT[0].t4 VDD.t812 VDD.t811 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3485 a_1533_n953.t25 WWLD[1].t20 a_1522_4445.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3486 a_3247_1457.t1 a_3152_1442.t3 VDD.t1796 VDD.t1795 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3487 a_8327_196.t0 WWL[14].t23 a_8595_4887.t19 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3488 a_2097_3425.t2 a_2002_3410.t3 VDD.t990 VDD.t989 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3489 a_7190_n953.t40 RWL[3].t12 a_7190_2943.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3490 a_7642_2662.t1 RWLB[4].t10 a_7190_n953.t35 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3491 a_7039_n5850.t0 PRE_CLSA.t93 VDD.t256 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3492 a_935_n1770.t2 a_1120_4887.t27 a_1128_n1770.t0 VSS.t2267 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3493 a_7067_4148.t0 VSS.t582 a_6615_n953.t15 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3494 a_1427_2647.t2 WWL[4].t20 a_1695_4887.t24 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3495 a_6122_n30.t2 a_6027_n45.t4 VDD.t1497 VDD.t1496 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3496 a_852_4133.t0 WWLD[2].t20 a_1120_4887.t20 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3497 a_3727_3169.t0 WWL[2].t20 a_3995_4887.t3 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3498 a_2002_2165.t2 WWL[6].t23 a_2270_4887.t21 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3499 VDD.t734 a_1522_n30.t4 a_1427_n45.t0 VDD.t733 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3500 VSS.t1025 a_n2677_n4378.t7 a_n2677_n5092.t1 VSS.t1019 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3501 a_8915_n953.t25 RWL[4].t13 a_8915_2662.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3502 a_6040_n953.t44 RWL[6].t7 a_6040_2180.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3503 a_5917_975.t0 RWLB[11].t14 a_5465_n953.t23 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3504 a_4675_n8583.t0 PRE_CLSA.t94 VDD.t258 VDD.t257 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3505 VSS.t1082 a_3231_n4378.t0 a_3231_n4378.t1 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3506 SA_OUT[4].t1 a_2610_n1371.t4 a_2853_n1770.t0 VSS.t1122 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3507 a_6697_n1053.t1 a_6602_n1068.t4 VDD.t1685 VDD.t1684 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3508 VSS.t1556 a_1522_2421.t5 a_1427_2406.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3509 a_1440_1216.t1 a_1427_1201.t5 VSS.t1532 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3510 VSS.t2008 a_3822_2943.t4 a_3727_2928.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3511 a_7847_n30.t0 a_7752_n45.t4 VDD.t794 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3512 VDD.t260 PRE_CLSA.t95 ADC9_OUT[0].t0 VDD.t259 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3513 a_2893_n2086.t1 a_2652_n2234.t4 VSS.t1174 VSS.t1173 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3514 a_8217_2421.t0 RWLB[5].t11 a_7765_n953.t23 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3515 a_13934_n5338.t0 SAEN.t83 a_14131_n5293.t0 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3516 a_11984_n5338.t1 Iref1.t8 a_12043_n5293.t1 VSS.t2227 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3517 VSS.t1467 a_947_4148.t3 a_1317_4148.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3518 VSS.t1768 a_2097_2180.t3 a_2467_2180.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3519 VDD.t962 a_6122_4445.t4 a_6027_4430.t1 VDD.t961 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3520 a_6122_975.t1 a_6027_960.t5 VSS.t2527 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3521 a_8217_n271.t0 VSS.t581 a_7765_n953.t9 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3522 a_8792_n812.t0 VSS.t580 a_8340_n953.t20 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3523 VSS.t1125 a_5547_2662.t5 a_5452_2647.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3524 a_2577_n827.t0 WWLD[6].t23 a_2845_4887.t6 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3525 VSS.t409 a_7847_3184.t5 a_7752_3169.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3526 a_5630_n6503.t1 a_5743_n6391# a_5595_n6849.t1 VSS.t207 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3527 VSS.t1923 a_n314_n4378.t1 a_n314_n4378.t2 VSS.t1922 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3528 a_5465_1939.t0 a_5452_1924.t5 VSS.t1176 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3529 a_2672_1698.t2 a_2577_1683.t4 VSS.t2105 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3530 a_9008_n953.t1 WWLD[5].t25 a_8997_n512.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3531 a_1522_3666.t0 a_1427_3651.t4 VSS.t1269 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3532 a_6697_1457.t1 a_6602_1442.t3 VDD.t1558 VDD.t1557 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3533 VDD.t738 a_8997_693.t5 a_8902_678.t1 VDD.t737 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3534 a_11776_n7216.t1 ADC13_OUT[2].t3 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3535 SA_OUT[2].t2 a_1460_n1371.t4 VDD.t2259 VDD.t2258 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3536 a_1317_3907.t0 VSS.t579 a_865_n953.t12 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3537 VDD.t1908 a_2672_2943.t5 a_2577_2928.t1 VDD.t1907 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3538 a_1337_n5338.t1 Iref1.t9 a_1396_n5293.t1 VSS.t2228 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3539 a_5452_2165.t0 WWL[6].t24 a_5720_4887.t23 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3540 a_1892_n30.t1 RWLB[15].t10 a_1440_n953.t32 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3541 a_3617_2943.t1 RWLB[3].t8 a_3165_n953.t37 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3542 a_14072_n7203.t1 Iref2.t6 a_14131_n6847.t1 VSS.t1984 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3543 a_5768_n2086.t1 a_5527_n2234.t4 VSS.t1764 VSS.t1763 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3544 a_742_2180.t0 RWLB[6].t9 a_290_n953.t41 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3545 VSS.t836 a_1522_1939.t4 a_1892_1939.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3546 a_2002_437.t2 WWL[13].t21 a_2270_4887.t26 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3547 a_7765_n953.t48 RWL[13].t10 a_7765_452.t1 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3548 VDD.t2276 a_n1233_n7216.t3 ADC2_OUT[2].t1 VDD.t1590 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3549 a_2085_n1770.t2 a_2270_4887.t27 a_2278_n1770.t1 VSS.t2423 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3550 a_6133_n953.t19 WWLD[0].t22 a_6122_4686.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3551 a_7765_3666.t1 a_7752_3651.t5 VSS.t1841 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3552 a_3247_1457.t0 a_3152_1442.t4 VSS.t2045 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3553 VSS.t2323 a_6697_452.t4 a_6602_437.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3554 VSS.t1159 a_6268_n2426.t7 a_7959_n7825.t1 VSS.t1156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3555 a_9405_n8583.t2 ADC11_OUT[3].t4 a_9475_n8071.t1 VSS.t2091 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3556 VSS.t1736 a_7272_2943.t5 a_7177_2928.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3557 VDD.t1407 a_1522_2662.t4 a_1427_2647.t1 VDD.t1406 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3558 VSS.t1329 a_5547_2180.t3 a_5917_2180.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3559 a_372_1698.t2 a_277_1683.t4 VDD.t1876 VDD.t1875 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3560 a_8915_n953.t0 RWL[15].t9 a_8915_n30.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3561 VSS.t2135 a_7418_n2426.t7 a_10327_n7825.t1 VSS.t2132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3562 a_2015_4686.t1 a_2002_4671.t4 VSS.t1810 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3563 a_1892_1698.t0 RWLB[8].t11 a_1440_n953.t29 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3564 a_3258_n953.t18 WWL[14].t24 a_3247_211.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3565 a_n2415_n7216.t2 ADC1_OUT[2].t4 a_n2345_n7203.t2 VSS.t1661 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3566 a_7994_n8026.t1 VCLP.t80 a_7959_n7825.t0 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3567 a_8915_1939.t0 a_8902_1924.t3 VSS.t1473 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3568 a_290_693.t1 a_277_678.t5 VSS.t2259 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3569 a_3247_4686.t2 a_3152_4671.t3 VDD.t1845 VDD.t1844 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3570 VSS.t1745 a_6122_2662.t5 a_6027_2647.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3571 a_6040_1457.t0 a_6027_1442.t5 VSS.t1583 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3572 a_2672_1216.t2 a_2577_1201.t4 VSS.t1765 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3573 a_5547_211.t0 a_5452_196.t5 VSS.t159 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3574 VDD.t1597 a_n2415_n4483.t4 ADC1_OUT[0].t2 VDD.t1596 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3575 a_4983_n953.t17 WWL[14].t25 a_4972_211.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3576 a_290_2943.t0 a_277_2928.t5 VSS.t769 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3577 a_1317_3425.t1 RWLB[1].t7 a_865_n953.t3 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3578 VSS.t903 a_2672_2421.t5 a_3042_2421.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3579 a_2467_1457.t0 RWLB[9].t11 a_2015_n953.t28 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3580 VSS.t362 SAEN.t84 a_n279_n3770.t0 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3581 a_4877_4133.t0 WWLD[2].t21 a_5145_4887.t11 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3582 a_4315_693.t1 a_4302_678.t5 VSS.t2290 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3583 a_1522_n30.t1 a_1427_n45.t4 VDD.t1099 VDD.t1098 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3584 a_1129_n4483.t0 PRE_CLSA.t96 VDD.t262 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3585 a_1440_4445.t1 a_1427_4430.t5 VSS.t1128 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3586 a_4192_2943.t0 RWLB[3].t9 a_3740_n953.t33 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3587 a_12736_n8026.t2 a_12963_n8583.t4 ADC14_OUT[3].t2 VSS.t1538 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3588 a_3165_n953.t3 VSS.t578 a_3165_3907.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3589 a_6122_3907.t0 a_6027_3892.t4 VSS.t1342 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3590 a_9475_n4470.t0 SAEN.t85 a_9672_n4114.t0 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3591 a_277_3169.t0 WWL[2].t21 a_545_4887.t25 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3592 a_6918_n2086.t0 a_6677_n2234.t4 VSS.t2069 VSS.t2068 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3593 VDD.t1187 a_947_4148.t4 a_852_4133.t1 VDD.t1186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3594 VDD.t522 a_7272_3184.t4 a_7177_3169.t1 VDD.t521 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3595 a_8422_2943.t1 a_8327_2928.t4 VSS.t2094 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3596 VDD.t1513 a_2097_2180.t4 a_2002_2165.t0 VDD.t1512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3597 a_6697_1939.t1 a_6602_1924.t5 VSS.t1382 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3598 a_6040_211.t0 a_6027_196.t5 VSS.t1152 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3599 a_3727_437.t2 WWL[13].t22 a_3995_4887.t20 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3600 a_3266_n3770.t2 a_3493_n4483.t3 ADC6_OUT[0].t1 VSS.t461 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3601 a_947_2943.t1 a_852_2928.t4 VSS.t1284 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3602 VSS.t1958 a_6122_2180.t4 a_6492_2180.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3603 a_7752_n827.t0 WWLD[6].t24 a_8020_4887.t6 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3604 VSS.t1956 a_4972_4148.t4 a_5342_4148.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3605 a_2108_n953.t21 WWL[4].t21 a_2097_2662.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3606 a_6027_2406.t0 WWL[5].t19 a_6295_4887.t10 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3607 a_372_1216.t2 a_277_1201.t5 VDD.t323 VDD.t322 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3608 a_1522_975.t1 a_1427_960.t5 VSS.t997 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3609 a_6697_4686.t1 a_6602_4671.t3 VDD.t994 VDD.t993 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3610 VSS.t1018 a_372_3184.t4 a_742_3184.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3611 a_1892_1216.t1 RWLB[10].t11 a_1440_n953.t36 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3612 a_7272_452.t1 a_7177_437.t5 VSS.t467 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3613 a_6027_n286.t2 WWLD[4].t18 a_6295_4887.t13 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3614 VSS.t2026 a_8997_4148.t5 a_8902_4133.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3615 a_10659_n7203.t0 a_5632_n6430# a_10856_n6847.t0 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3616 a_2590_n953.t0 RWL[0].t14 a_2590_3666.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3617 a_8997_3666.t0 a_8902_3651.t4 VSS.t1217 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3618 VSS.t252 a_3822_693.t5 a_3727_678.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3619 VDD.t2104 a_4397_693.t5 a_4302_678.t2 VDD.t2103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3620 a_5342_3907.t0 VSS.t577 a_4890_n953.t9 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3621 VDD.t610 a_6697_2943.t4 a_6602_2928.t1 VDD.t609 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3622 a_5917_1457.t1 RWLB[9].t12 a_5465_n953.t32 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3623 VDD.t900 a_372_n30.t4 a_277_n45.t0 VDD.t899 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3624 a_4675_n5850.t2 ADC7_OUT[1].t4 a_4745_n5338.t2 VSS.t1262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3625 a_n52_n5850.t2 ADC3_OUT[1].t4 a_18_n5338.t2 VSS.t1123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3626 VDD.t1220 PRE_A.t13 a_7843_n2422.t2 VDD.t1219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3627 VSS.t1809 a_6697_1939.t5 a_7067_1939.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3628 a_1129_n7216.t2 ADC4_OUT[2].t4 a_1199_n7203.t2 VSS.t1046 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3629 a_8327_4133.t0 WWLD[2].t22 a_8595_4887.t13 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3630 a_3165_n953.t9 VSS.t576 a_3165_n271.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3631 a_3247_4686.t1 a_3152_4671.t4 VSS.t1407 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3632 a_6615_n953.t4 VSS.t575 a_6615_3907.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3633 a_7642_2943.t0 RWLB[3].t10 a_7190_n953.t31 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3634 a_1427_2928.t0 WWL[3].t20 a_1695_4887.t0 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3635 a_4315_n953.t23 RWL[11].t7 a_4315_975.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3636 a_1533_n953.t12 WWL[5].t20 a_1522_2421.t0 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3637 VDD.t970 a_5547_2180.t4 a_5452_2165.t1 VDD.t969 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3638 VSS.t149 a_5547_693.t5 a_5917_693.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3639 a_7272_1457.t1 a_7177_1442.t4 VSS.t507 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3640 a_n3495_n5338.t0 SAEN.t86 a_n3298_n5293.t0 VSS.t336 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3641 a_3165_n953.t20 RWL[1].t10 a_3165_3425.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3642 a_6122_3425.t1 a_6027_3410.t4 VSS.t2087 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3643 a_9613_n8071.t0 VCLP.t81 a_9475_n8071.t2 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3644 a_7765_n953.t3 VSS.t574 a_7765_n1053.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3645 a_11776_n7216.t0 PRE_CLSA.t97 VDD.t263 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3646 a_7067_1698.t1 RWLB[8].t12 a_6615_n953.t34 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3647 a_852_1683.t0 WWL[8].t20 a_1120_4887.t19 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3648 VSS.t152 a_7272_211.t5 a_7642_211.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3649 a_6040_4686.t1 a_6027_4671.t5 VSS.t1048 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3650 a_11984_n5338.t0 VCLP.t82 a_11846_n5338.t1 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3651 a_5630_n3770.t1 VCLP.t83 a_5595_n4116.t0 VSS.t186 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3652 VSS.t2369 a_3247_3907.t5 a_3152_3892.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3653 a_8429_n8071.t1 Iref3.t15 a_8488_n8026.t1 VSS.t1979 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3654 a_9027_n1770.t0 SA_OUT[15].t4 a_8935_n1371.t2 VSS.t2084 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3655 a_4983_n953.t25 WWL[6].t25 a_4972_2180.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3656 VSS.t1539 a_947_975.t5 a_852_960.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3657 VDD.t724 a_2311_n8583.t4 ADC5_OUT[3].t1 VDD.t723 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3658 a_n3792_n5293.t2 a_n3565_n5850.t4 ADC0_OUT[1].t1 VSS.t427 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3659 a_2672_4445.t0 a_2577_4430.t4 VSS.t1111 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3660 a_3833_n953.t16 WWLD[2].t23 a_3822_4148.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3661 VDD.t2069 PRE_SRAM.t33 a_383_n953.t3 VDD.t2068 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3662 a_2467_4686.t0 VSS.t573 a_2015_n953.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3663 VDD.t1230 a_6122_2421.t4 a_6027_2406.t2 VDD.t1229 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3664 a_4877_n45.t2 WWL[15].t23 a_5145_4887.t9 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3665 a_13637_n6503.t0 a_13864_n7216.t4 ADC15_OUT[2].t2 VSS.t1409 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3666 VSS.t2430 a_4397_n1053.t5 a_4302_n1068.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3667 VSS.t1593 a_947_1698.t3 a_1317_1698.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3668 a_n3357_n7203.t1 Iref2.t7 a_n3298_n6847.t1 VSS.t824 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3669 a_n2345_n8071.t0 SAEN.t87 a_n2148_n8026.t0 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3670 a_n1460_n5293.t1 VCLP.t84 a_n1495_n5092.t0 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3671 a_13033_n7203.t0 a_5632_n6430# a_13230_n6847.t0 VSS.t348 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3672 a_4192_693.t0 RWLB[12].t9 a_3740_n953.t23 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3673 a_6615_n953.t3 VSS.t572 a_6615_n271.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3674 a_10362_n6503.t2 a_5743_n6391# a_10327_n6849.t1 VSS.t210 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3675 a_5342_3425.t0 RWLB[1].t8 a_4890_n953.t33 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3676 a_6492_1457.t1 RWLB[9].t13 a_6040_n953.t32 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3677 a_3701_n5338.t1 Iref1.t10 a_3760_n5293.t1 VSS.t2229 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3678 a_13864_n4483.t2 ADC15_OUT[0].t4 VDD.t1031 VDD.t1030 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3679 VSS.t1757 a_947_n812.t3 a_1317_n812.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3680 a_5558_n953.t14 WWL[7].t24 a_5547_1939.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3681 a_7190_n953.t8 VSS.t571 a_7190_3907.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3682 VSS.t2243 a_2672_3666.t4 a_2577_3651.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3683 a_7765_n953.t19 RWL[9].t13 a_7765_1457.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3684 a_6615_n953.t21 RWL[1].t11 a_6615_3425.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3685 VDD.t1668 a_8422_4148.t4 a_8327_4133.t2 VDD.t1667 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3686 a_372_4445.t1 a_277_4430.t5 VDD.t1984 VDD.t1983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3687 a_1440_211.t1 a_1427_196.t5 VSS.t1895 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 a_6065_n5338.t1 Iref1.t11 a_6124_n5293.t1 VSS.t2230 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3689 VSS.t2294 a_3247_n271.t5 a_3152_n286.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3690 a_1892_4445.t0 VSS.t570 a_1440_n953.t2 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3691 VSS.t1395 a_8993_n2422.t1 a_8993_n2422.t2 VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3692 a_n2415_n4483.t1 ADC1_OUT[0].t3 a_n2345_n4470.t2 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3693 a_3822_n812.t1 a_3727_n827.t5 VDD.t1986 VDD.t1985 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3694 a_7067_1216.t1 RWLB[10].t12 a_6615_n953.t41 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3695 VSS.t1213 a_5543_n2422.t7 a_6777_n5092.t1 VSS.t1207 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3696 a_6133_n953.t11 WWL[4].t22 a_6122_2662.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3697 a_852_1201.t0 WWL[10].t21 a_1120_4887.t5 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3698 VSS.t938 a_475_n2132.t2 a_453_n2086.t0 VSS.t937 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3699 a_277_960.t0 WWL[11].t25 a_545_4887.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3700 VSS.t2447 a_3822_3907.t4 a_3727_3892.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3701 VSS.t2449 a_3247_3425.t5 a_3152_3410.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3702 VSS.t1842 a_4397_1457.t5 a_4302_1442.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3703 a_2672_452.t0 a_2577_437.t5 VSS.t1975 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3704 a_5857_n7216.t2 ADC8_OUT[2].t3 VDD.t472 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3705 a_5917_4686.t0 VSS.t569 a_5465_n953.t2 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3706 a_8217_n30.t0 RWLB[15].t11 a_7765_n953.t41 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3707 a_2015_2662.t0 a_2002_2647.t4 VSS.t410 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3708 VSS.t2507 a_3227_n2234.t4 a_3350_n2132.t0 VSS.t2506 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3709 VDD.t264 PRE_CLSA.t98 ADC4_OUT[2].t0 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3710 a_2077_n2234.t1 Din[3].t1 VSS.t1423 VSS.t1422 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3711 VSS.t1866 a_947_1216.t3 a_1317_1216.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3712 a_6602_3892.t2 WWLD[3].t23 a_6870_4887.t9 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3713 a_3247_2662.t2 a_3152_2647.t3 VDD.t1471 VDD.t1470 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3714 a_7190_n953.t4 VSS.t568 a_7190_n271.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3715 a_7272_4686.t2 a_7177_4671.t4 VSS.t1487 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3716 VDD.t266 PRE_CLSA.t99 ADC5_OUT[3].t2 VDD.t265 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3717 a_8340_n953.t26 RWL[11].t8 a_8340_975.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3718 VSS.t2241 a_947_211.t5 a_1317_211.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3719 VSS.t2213 a_3822_n30.t5 a_3727_n45.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3720 VDD.t1662 a_2672_3907.t5 a_2577_3892.t2 VDD.t1661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3721 a_2672_n512.t2 a_2577_n527.t5 VDD.t1934 VDD.t1933 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3722 a_7190_n953.t23 RWL[1].t12 a_7190_3425.t1 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3723 SA_OUT[2].t0 PRE_VLSA.t41 VDD.t1109 VDD.t1108 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3724 a_865_n953.t25 RWL[11].t9 a_865_975.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3725 a_7847_975.t1 a_7752_960.t5 VSS.t2520 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3726 a_11846_n5338.t0 SAEN.t88 a_12043_n5293.t0 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3727 a_3165_n812.t1 a_3152_n827.t5 VSS.t959 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3728 a_383_n953.t18 WWL[3].t21 a_372_2943.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3729 a_1440_2421.t1 a_1427_2406.t5 VSS.t1350 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3730 a_5547_693.t1 a_5452_678.t4 VDD.t2100 VDD.t2099 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3731 a_290_n953.t35 EN.t10 a_n3827_n4378.t3 VSS.t1950 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3732 VSS.t866 a_6102_n2234.t4 a_6225_n2132.t0 VSS.t865 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3733 VDD.t2199 a_3822_n1053.t5 a_3727_n1068.t2 VDD.t2198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3734 a_3822_3184.t2 a_3727_3169.t4 VSS.t2003 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3735 VSS.t2298 a_4397_975.t3 a_4767_975.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3736 a_3727_3651.t2 WWL[0].t22 a_3995_4887.t26 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3737 a_4877_1683.t2 WWL[8].t21 a_5145_4887.t10 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3738 a_1440_n271.t1 a_1427_n286.t5 VSS.t2090 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3739 VSS.t1685 a_3822_n271.t4 a_3727_n286.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3740 a_9008_n953.t14 WWLD[2].t24 a_8997_4148.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3741 VSS.t2461 a_7272_3907.t5 a_7177_3892.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3742 VSS.t2100 a_8568_n2426.t6 a_12701_n4116.t1 VSS.t2095 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3743 a_10659_n4470.t0 SAEN.t89 a_10856_n4114.t0 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3744 a_7752_n1068.t0 WWLD[7].t20 a_8020_4887.t22 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3745 VSS.t2001 a_4972_975.t5 a_4877_960.t2 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3746 VDD.t1342 a_947_1698.t4 a_852_1683.t1 VDD.t1341 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3747 VSS.t2495 a_3822_3425.t4 a_3727_3410.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3748 a_2097_n30.t2 a_2002_n45.t5 VSS.t1363 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3749 a_1199_n5338.t0 SAEN.t90 a_1396_n5293.t0 VSS.t342 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3750 VSS.t1917 a_8422_n1053.t5 a_8327_n1068.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3751 VSS.t383 a_3247_n512.t4 a_3617_n512.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3752 a_6492_4686.t0 VSS.t567 a_6040_n953.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3753 a_8340_975.t1 a_8327_960.t5 VSS.t2184 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3754 a_1129_n4483.t1 ADC4_OUT[0].t3 a_1199_n4470.t2 VSS.t1638 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3755 a_6697_2662.t1 a_6602_2647.t4 VDD.t1944 VDD.t1943 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3756 a_4890_2180.t0 a_4877_2165.t5 VSS.t1941 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3757 VSS.t1 a_4972_1698.t5 a_5342_1698.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 VDD.t1501 a_947_n812.t4 a_852_n827.t1 VDD.t1500 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3759 a_3740_4148.t1 a_3727_4133.t5 VSS.t1070 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3760 a_6122_4148.t1 a_6027_4133.t5 VDD.t2247 VDD.t2246 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3761 a_7272_2180.t1 a_7177_2165.t5 VDD.t2225 VDD.t2224 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3762 VSS.t1529 a_2672_452.t5 a_3042_452.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3763 a_11984_n7203.t1 Iref2.t8 a_12043_n6847.t1 VSS.t825 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3764 VSS.t1537 a_4377_n2234.t4 a_4500_n2132.t0 VSS.t1536 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3765 a_7765_n953.t5 VSS.t566 a_7765_4686.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3766 a_8997_3184.t2 a_8902_3169.t5 VDD.t864 VDD.t863 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3767 VSS.t1850 a_7847_3666.t5 a_7752_3651.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3768 VSS.t2142 a_8997_1698.t5 a_8902_1683.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3769 VDD.t814 a_2672_n271.t5 a_2577_n286.t2 VDD.t813 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3770 a_6602_3410.t0 WWL[1].t24 a_6870_4887.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3771 a_3227_n2234.t1 Din[5].t1 VSS.t1235 VSS.t1234 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3772 VSS.t111 a_4972_n812.t5 a_5342_n812.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3773 VDD.t520 a_3822_1457.t5 a_3727_1442.t1 VDD.t519 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3774 VSS.t2205 a_8997_n812.t5 a_8902_n827.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3775 a_6615_n812.t1 a_6602_n827.t4 VSS.t1616 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3776 a_7067_4445.t0 VSS.t565 a_6615_n953.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3777 VDD.t1660 a_2672_3425.t5 a_2577_3410.t2 VDD.t1659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3778 a_3247_2662.t1 a_3152_2647.t4 VSS.t1717 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3779 a_1603_n2086.t1 WE.t24 a_1533_n953.t15 VSS.t2397 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3780 a_852_4430.t2 WWLD[1].t21 a_1120_4887.t21 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3781 a_8327_1683.t0 WWL[8].t22 a_8595_4887.t12 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3782 VSS.t2350 a_7272_n271.t5 a_7177_n286.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3783 a_1337_n7203.t1 Iref2.t9 a_1396_n6847.t1 VSS.t826 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3784 a_7847_n812.t1 a_7752_n827.t3 VDD.t767 VDD.t766 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3785 VSS.t1351 a_4397_4686.t5 a_4302_4671.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3786 a_2845_4887.t20 PRE_SRAM.t34 VDD.t2071 VDD.t2070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3787 a_4877_1201.t0 WWL[10].t22 a_5145_4887.t3 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3788 VSS.t237 a_8422_n30.t4 a_8792_n30.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3789 a_13864_n4483.t0 PRE_CLSA.t100 VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3790 VSS.t1501 a_7252_n2234.t3 a_7375_n2132.t0 VSS.t1500 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3791 VSS.t1429 a_8422_1457.t5 a_8327_1442.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3792 a_10797_n8071.t0 VCLP.t85 a_10659_n8071.t1 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3793 a_13637_n3770.t2 a_13864_n4483.t3 ADC15_OUT[0].t1 VSS.t1236 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3794 a_4408_n953.t25 WWLD[7].t21 a_4397_n1053.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3795 VSS.t479 a_7272_3425.t5 a_7177_3410.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3796 a_290_n953.t9 VSS.t564 a_290_n512.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3797 VDD.t1097 a_4675_n8583.t4 ADC7_OUT[3].t2 VDD.t1096 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3798 VSS.t63 a_947_4445.t4 a_1317_4445.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3799 a_6040_2662.t1 a_6027_2647.t5 VSS.t1558 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3800 VDD.t1628 a_947_1216.t4 a_852_1201.t2 VDD.t1627 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3801 a_3617_n30.t0 RWLB[15].t12 a_3165_n953.t34 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3802 a_13033_n4470.t0 SAEN.t91 a_13230_n4114.t0 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3803 a_10362_n3770.t1 VCLP.t86 a_10327_n4116.t0 VSS.t190 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3804 VSS.t2362 a_3822_n512.t5 a_4192_n512.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3805 a_4478_n2086.t0 WE.t25 a_4408_n953.t8 VSS.t2398 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3806 a_4397_n812.t2 a_4302_n827.t5 VSS.t2253 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3807 a_2672_2421.t1 a_2577_2406.t4 VSS.t931 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3808 a_8902_1924.t2 WWL[7].t25 a_9170_4887.t8 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 VSS.t56 a_4972_1216.t5 a_5342_1216.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3810 a_958_n953.t6 WWL[12].t22 a_947_693.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3811 a_3833_n953.t23 WWL[8].t23 a_3822_1698.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3812 a_2672_n271.t1 a_2577_n286.t4 VSS.t1195 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3813 a_5465_n512.t1 a_5452_n527.t5 VSS.t2139 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3814 a_2467_2662.t1 RWLB[4].t11 a_2015_n953.t36 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3815 VSS.t2061 a_8997_1216.t5 a_8902_1201.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3816 a_7765_211.t1 a_7752_196.t5 VSS.t1332 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3817 VSS.t1579 a_867_n4378.t7 a_867_n5092.t1 VSS.t1573 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3818 VDD.t2140 a_6697_3907.t4 a_6602_3892.t1 VDD.t2139 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3819 a_5452_437.t2 WWL[13].t23 a_5720_4887.t14 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3820 VDD.t335 a_7827_n2234.t4 a_7950_n2132.t1 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3821 VDD.t2122 a_4397_975.t4 a_4302_960.t2 VDD.t2121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3822 a_5857_n7216.t0 PRE_CLSA.t101 VDD.t269 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3823 a_3833_n953.t1 WWLD[6].t25 a_3822_n812.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3824 a_947_211.t1 a_852_196.t4 VDD.t930 VDD.t929 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3825 VSS.t367 SAEN.t92 a_n1460_n6503.t0 VSS.t350 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3826 a_7190_n812.t1 a_7177_n827.t5 VSS.t1720 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3827 a_4972_4148.t1 a_4877_4133.t3 VSS.t1911 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3828 a_4890_n953.t29 RWL[2].t14 a_4890_3184.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3829 a_8327_1201.t0 WWL[10].t23 a_8595_4887.t3 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3830 VSS.t2189 a_8422_975.t5 a_8792_975.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3831 a_8997_452.t1 a_8902_437.t5 VSS.t842 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3832 a_n3565_n8583.t2 ADC0_OUT[3].t4 VDD.t916 VDD.t915 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3833 a_2753_n2086.t0 WE.t26 a_2683_n953.t7 VSS.t2399 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3834 a_4408_n953.t14 WWL[9].t23 a_4397_1457.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3835 a_2015_975.t1 a_2002_960.t5 VSS.t880 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3836 a_372_2421.t2 a_277_2406.t5 VDD.t680 VDD.t679 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3837 VDD.t892 a_6122_211.t5 a_6027_196.t1 VDD.t891 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3838 VDD.t313 a_3247_n512.t5 a_3152_n527.t2 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3839 a_277_3651.t2 WWL[0].t23 a_545_4887.t20 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3840 VDD.t1916 a_8422_1698.t5 a_8327_1683.t2 VDD.t1915 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3841 VDD.t2146 a_7272_3666.t5 a_7177_3651.t2 VDD.t2145 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3842 a_1892_2421.t0 RWLB[5].t12 a_1440_n953.t41 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3843 a_6708_n953.t9 WWL[14].t26 a_6697_211.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3844 a_372_n271.t1 a_277_n286.t5 VDD.t2281 VDD.t2280 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3845 a_8429_n5338.t0 VCLP.t87 a_8291_n5338.t1 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3846 a_742_n1053.t0 VSS.t563 a_290_n953.t5 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3847 VSS.t2160 a_7272_n512.t5 a_7642_n512.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3848 VSS.t2477 a_8997_n30.t5 a_9367_n30.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3849 a_1892_n271.t0 VSS.t562 a_1440_n953.t4 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3850 a_13171_n8071.t0 VCLP.t88 a_13033_n8071.t1 VSS.t222 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3851 a_7847_n812.t2 a_7752_n827.t4 VSS.t1139 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3852 a_2015_2943.t0 a_2002_2928.t4 VSS.t2027 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3853 a_3740_975.t1 a_3727_960.t5 VSS.t2372 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3854 a_947_3907.t2 a_852_3892.t3 VDD.t534 VDD.t533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3855 VSS.t1756 a_1522_3184.t5 a_1427_3169.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3856 a_1522_1457.t1 a_1427_1442.t5 VDD.t832 VDD.t831 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3857 a_4890_n953.t0 RWL[15].t10 a_4890_n30.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3858 VDD.t1958 a_8422_n812.t5 a_8327_n827.t2 VDD.t1957 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3859 a_8915_n512.t1 a_8902_n527.t3 VSS.t1688 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3860 a_5465_n953.t18 RWL[3].t13 a_5465_2943.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3861 a_5917_2662.t0 RWLB[4].t12 a_5465_n953.t39 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3862 a_10589_n7216.t2 ADC12_OUT[2].t3 VDD.t1277 VDD.t1276 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3863 VSS.t2207 a_372_3666.t5 a_742_3666.t1 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3864 a_3042_2180.t0 RWLB[6].t10 a_2590_n953.t40 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3865 VDD.t45 a_6697_n271.t5 a_6602_n286.t1 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3866 a_2683_n953.t2 WWLD[5].t26 a_2672_n512.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3867 VDD.t1027 a_3822_4686.t5 a_3727_4671.t2 VDD.t1026 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3868 a_8217_3184.t1 RWLB[2].t12 a_7765_n953.t40 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3869 a_3247_2943.t2 a_3152_2928.t3 VDD.t1570 VDD.t1569 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3870 VSS.t2322 a_372_n512.t5 a_277_n527.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3871 a_3833_n953.t8 WWL[10].t24 a_3822_1216.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3872 a_5628_n2086.t0 WE.t27 a_5558_n953.t12 VSS.t2410 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3873 a_4315_n953.t41 RWL[6].t8 a_4315_2180.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3874 SA_OUT[0].t1 a_310_n1371.t4 VDD.t1183 VDD.t1182 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3875 VDD.t25 a_6697_3425.t5 a_6602_3410.t2 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3876 a_7272_2662.t1 a_7177_2647.t4 VSS.t1255 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3877 VDD.t2166 a_8977_n2234.t4 a_9100_n2132.t1 VDD.t2165 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3878 a_4877_4430.t0 WWLD[1].t22 a_5145_4887.t15 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3879 VSS.t1233 a_2097_2943.t5 a_2002_2928.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3880 a_n2415_n4483.t0 PRE_CLSA.t102 VDD.t271 VDD.t270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3881 VSS.t1170 a_8422_4686.t5 a_8327_4671.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3882 a_865_n953.t38 RWL[13].t11 a_865_452.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3883 a_8433_n953.t16 WWL[13].t24 a_8422_452.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3884 VDD.t1222 PRE_A.t14 a_n3827_n4378.t2 VDD.t1221 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3885 a_6870_4887.t3 PRE_SRAM.t35 VDD.t2073 VDD.t2072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3886 VDD.t17 a_947_4445.t5 a_852_4430.t1 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3887 a_6697_n512.t2 a_6602_n527.t5 VSS.t2510 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3888 a_6602_n45.t2 WWL[15].t24 a_6870_4887.t24 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3889 a_8433_n953.t19 WWLD[7].t22 a_8422_n1053.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3890 VSS.t2144 a_947_2180.t5 a_852_2165.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3891 VSS.t843 a_8997_452.t5 a_9367_452.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3892 VSS.t2426 a_4972_4445.t5 a_5342_4445.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3893 VDD.t1996 a_8422_1216.t5 a_8327_1201.t2 VDD.t1995 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3894 a_958_n953.t24 WWLD[7].t23 a_947_n1053.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3895 a_4397_3907.t1 a_4302_3892.t4 VDD.t838 VDD.t837 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3896 a_8915_n953.t17 RWL[3].t14 a_8915_2943.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3897 a_3740_n953.t29 RWL[7].t13 a_3740_1939.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3898 a_8340_n953.t41 RWL[12].t11 a_8340_693.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3899 VSS.t2434 a_n1495_n4378.t0 a_n1495_n4378.t1 VSS.t2433 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3900 a_9008_n953.t15 WWL[8].t24 a_8997_1698.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3901 VDD.t972 a_7847_211.t5 a_7752_196.t0 VDD.t971 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3902 a_3563_n5338.t0 SAEN.t93 a_3760_n5293.t0 VSS.t346 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3903 VSS.t1231 a_8997_4445.t5 a_8902_4430.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3904 VSS.t93 a_n3827_n4378.t6 a_n3827_n6849.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3905 a_1120_4887.t26 PRE_SRAM.t36 a_958_n953.t22 VDD.t2074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3906 a_6697_2943.t2 a_6602_2928.t4 VDD.t1191 VDD.t1190 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3907 VSS.t1734 a_7272_693.t4 a_7177_678.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3908 VDD.t272 PRE_CLSA.t103 ADC14_OUT[1].t0 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3909 a_947_3425.t2 a_852_3410.t3 VDD.t598 VDD.t597 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3910 a_6492_2662.t1 RWLB[4].t13 a_6040_n953.t39 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3911 VSS.t102 a_4393_n2422.t6 a_4413_n6849.t1 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3912 a_9008_n953.t9 WWLD[6].t26 a_8997_n812.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3913 a_5465_n953.t1 RWL[15].t11 a_5465_n30.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3914 a_5927_n5338.t0 SAEN.t94 a_6124_n5293.t0 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3915 a_7765_n953.t28 RWL[4].t14 a_7765_2662.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3916 a_4408_n953.t21 WWLD[0].t23 a_4397_4686.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3917 a_8327_4430.t2 WWLD[1].t23 a_8595_4887.t17 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3918 a_3740_1698.t0 a_3727_1683.t5 VSS.t1985 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3919 a_6122_1698.t2 a_6027_1683.t5 VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3920 a_11549_n8026.t2 a_11776_n8583.t4 ADC13_OUT[3].t2 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3921 VSS.t926 a_5547_2943.t5 a_5452_2928.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3922 VSS.t2313 a_7843_n2422.t0 a_7843_n2422.t1 VSS.t2312 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3923 a_n3357_n8071.t0 VCLP.t89 a_n3495_n8071.t1 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3924 a_3247_2943.t1 a_3152_2928.t4 VSS.t871 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3925 a_372_2180.t1 a_277_2165.t4 VSS.t483 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3926 a_8433_n953.t20 WWL[9].t24 a_8422_1457.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3927 a_3701_n7203.t1 Iref2.t10 a_3760_n6847.t1 VSS.t827 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3928 a_14072_n7203.t0 a_5743_n6391# a_13934_n7203.t2 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3929 a_7067_2421.t0 RWLB[5].t13 a_6615_n953.t22 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3930 a_4675_n5850.t0 PRE_CLSA.t104 VDD.t273 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3931 a_n3565_n4483.t0 PRE_CLSA.t105 VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3932 VSS.t2022 a_2672_3184.t5 a_3042_3184.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3933 a_852_2406.t0 WWL[5].t21 a_1120_4887.t3 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3934 a_3165_452.t0 a_3152_437.t5 VSS.t2054 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3935 a_n1233_n8583.t2 ADC2_OUT[3].t4 a_n1163_n8071.t2 VSS.t1879 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3936 a_383_n953.t8 WWLD[3].t24 a_372_3907.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 a_958_n953.t12 WWL[9].t25 a_947_1457.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3938 VDD.t924 a_1522_211.t5 a_1427_196.t1 VDD.t923 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3939 a_6133_n953.t12 WWL[15].t25 a_6122_n30.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3940 a_7067_n271.t1 VSS.t561 a_6615_n953.t11 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3941 a_2084_n5293.t1 VCLP.t90 a_2049_n5092.t0 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X3942 a_n1025_n4470.t1 Iref0.t8 a_n966_n4114.t1 VSS.t2224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3943 a_1522_4686.t2 a_1427_4671.t5 VDD.t450 VDD.t449 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3944 VSS.t2032 a_4397_2662.t5 a_4302_2647.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3945 a_4315_1457.t0 a_4302_1442.t4 VSS.t941 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3946 a_852_n286.t0 WWLD[4].t19 a_1120_4887.t9 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3947 a_6065_n7203.t1 Iref2.t11 a_6124_n6847.t1 VSS.t828 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X3948 a_3165_n1053.t0 a_3152_n1068.t5 VSS.t2186 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3949 VSS.t1488 a_4972_n30.t4 a_5342_n30.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3950 a_977_n1770.t1 SA_OUT[1].t4 a_885_n1371.t2 VSS.t1938 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3951 a_6040_2943.t1 a_6027_2928.t5 VSS.t818 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3952 a_3833_n953.t25 WWLD[1].t24 a_3822_4445.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3953 a_4397_3425.t2 a_4302_3410.t4 VDD.t1542 VDD.t1541 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3954 a_5547_1457.t1 a_5452_1442.t3 VDD.t800 VDD.t799 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3955 a_8327_n45.t2 WWL[15].t26 a_8595_4887.t11 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3956 a_9008_n953.t2 WWL[10].t25 a_8997_1216.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3957 a_372_452.t1 a_277_437.t5 VSS.t444 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3958 a_4890_452.t0 a_4877_437.t5 VSS.t814 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3959 a_9367_4148.t0 VSS.t560 a_8915_n953.t6 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3960 VDD.t546 a_1522_2943.t5 a_1427_2928.t2 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3961 VSS.t2288 a_947_2421.t4 a_1317_2421.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3962 a_7642_693.t1 RWLB[12].t10 a_7190_n953.t21 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3963 a_2702_n1770.t1 a_2683_n953.t27 a_2660_n1770.t1 VSS.t2166 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3964 a_4302_2165.t2 WWL[6].t26 a_4570_4887.t12 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3965 a_7272_211.t0 a_7177_196.t4 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3966 a_2311_n8583.t2 ADC5_OUT[3].t4 VDD.t720 VDD.t719 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3967 a_3152_4133.t2 WWLD[2].t25 a_3420_4887.t16 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3968 a_6027_3169.t0 WWL[2].t22 a_6295_4887.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3969 a_2467_2943.t0 RWLB[3].t11 a_2015_n953.t32 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3970 a_2108_n953.t16 WWL[13].t25 a_2097_452.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3971 a_n1233_n7216.t0 PRE_CLSA.t106 VDD.t276 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3972 a_8977_n2234.t1 Din[15].t1 VSS.t1367 VSS.t1366 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3973 a_8340_n953.t43 RWL[6].t9 a_8340_2180.t1 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3974 VSS.t369 SAEN.t95 a_n1460_n3770.t0 VSS.t368 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X3975 a_1522_1939.t0 a_1427_1924.t4 VSS.t1805 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3976 a_865_n953.t43 RWL[6].t10 a_865_2180.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3977 a_2097_1457.t0 a_2002_1442.t5 VSS.t955 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3978 a_3740_1216.t0 a_3727_1201.t5 VSS.t1664 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3979 VDD.t1446 a_1129_n7216.t3 ADC4_OUT[2].t2 VDD.t1270 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X3980 VSS.t1921 a_6122_2943.t5 a_6027_2928.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3981 a_6122_1216.t2 a_6027_1201.t5 VDD.t808 VDD.t807 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3982 a_6040_n1053.t0 a_6027_n1068.t5 VSS.t1876 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3983 VSS.t853 a_4397_2180.t4 a_4767_2180.t0 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3984 a_3833_n953.t19 WWL[13].t26 a_3822_452.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3985 a_383_n953.t13 WWLD[4].t20 a_372_n271.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3986 VDD.t470 a_8422_4445.t5 a_8327_4430.t1 VDD.t469 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3987 VSS.t859 a_3247_4148.t4 a_3617_4148.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3988 a_2015_n953.t42 RWL[12].t12 a_2015_693.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3989 VSS.t1250 a_947_693.t4 a_852_678.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3990 VSS.t1943 a_4972_2180.t5 a_4877_2165.t0 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3991 VSS.t1771 a_5547_n30.t5 a_5452_n45.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3992 a_5577_n1770.t0 a_5558_n953.t27 a_5535_n1770.t0 VSS.t968 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3993 a_383_n953.t0 WWL[1].t25 a_372_3425.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3994 a_1533_n953.t3 WWL[2].t23 a_1522_3184.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3995 a_7765_1939.t1 a_7752_1924.t5 VSS.t1807 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3996 VSS.t437 a_4397_452.t5 a_4767_452.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3997 a_3822_3666.t1 a_3727_3651.t4 VSS.t1184 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3998 a_4972_1698.t1 a_4877_1683.t3 VSS.t249 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3999 a_3247_975.t2 a_3152_960.t4 VDD.t926 VDD.t925 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4000 VSS.t1901 a_372_211.t5 a_742_211.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4001 a_3740_n953.t43 RWL[12].t13 a_3740_693.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4002 a_3617_3907.t0 VSS.t559 a_3165_n953.t5 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4003 VDD.t586 a_3247_211.t5 a_3152_196.t0 VDD.t585 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4004 a_5145_4887.t20 PRE_SRAM.t37 a_4983_n953.t5 VDD.t2075 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4005 VSS.t2458 a_2049_n4378.t6 a_2049_n4116.t1 VSS.t2453 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4006 a_2127_n1770.t1 SA_OUT[3].t4 a_2035_n1371.t1 VSS.t1129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4007 a_4315_n1053.t1 a_4302_n1068.t5 VSS.t2445 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4008 VSS.t1131 a_2672_693.t4 a_2577_678.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4009 a_5917_2943.t1 RWLB[3].t12 a_5465_n953.t35 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4010 a_9178_n8026.t1 VCLP.t91 a_9143_n7825.t0 VSS.t223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4011 a_1440_n953.t1 RWL[15].t12 a_1440_n30.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4012 a_2108_n953.t18 WWL[3].t22 a_2097_2943.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4013 a_3852_n1770.t1 a_3833_n953.t27 a_3810_n1770.t2 VSS.t455 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4014 a_8433_n953.t8 WWLD[0].t24 a_8422_4686.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4015 a_8997_3666.t1 a_8902_3651.t5 VDD.t840 VDD.t839 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4016 a_5547_1457.t0 a_5452_1442.t4 VSS.t1167 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4017 VDD.t688 a_3822_2662.t5 a_3727_2647.t1 VDD.t687 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4018 a_8997_211.t1 a_8902_196.t5 VDD.t1390 VDD.t1389 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4019 a_n279_n8026.t2 a_n52_n8583.t4 ADC3_OUT[3].t1 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4020 VDD.t1248 a_6122_3184.t5 a_6027_3169.t2 VDD.t1247 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4021 a_7272_2943.t2 a_7177_2928.t4 VSS.t1137 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4022 a_958_n953.t20 WWLD[0].t25 a_947_4686.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4023 a_290_n953.t15 VSS.t558 a_290_4148.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4024 a_156_n5338.t1 Iref1.t12 a_215_n5293.t1 VSS.t2231 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4025 a_4315_4686.t1 a_4302_4671.t4 VSS.t1851 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4026 VSS.t1081 a_3822_4148.t5 a_4192_4148.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4027 a_8902_678.t2 WWL[12].t23 a_9170_4887.t6 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4028 a_4877_2406.t0 WWL[5].t22 a_5145_4887.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4029 VSS.t2112 a_8422_2662.t5 a_8327_2647.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4030 a_5547_4686.t1 a_5452_4671.t3 VDD.t1035 VDD.t1034 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4031 a_8340_1457.t1 a_8327_1442.t5 VSS.t1114 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4032 a_1317_693.t1 RWLB[12].t11 a_865_n953.t22 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4033 a_4877_n286.t2 WWLD[4].t21 a_5145_4887.t16 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4034 a_9008_n953.t18 WWLD[1].t25 a_8997_4445.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4035 a_290_3907.t1 a_277_3892.t5 VSS.t2329 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4036 VDD.t2114 a_947_2421.t5 a_852_2406.t2 VDD.t2113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4037 a_865_1457.t1 a_852_1442.t5 VSS.t2080 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4038 VSS.t988 a_6693_n2422.t7 a_9143_n5092.t1 VSS.t982 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4039 a_6727_n1770.t0 a_6708_n953.t27 a_6685_n1770.t2 VSS.t2305 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4040 a_4972_1216.t1 a_4877_1201.t3 VSS.t2359 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4041 a_5547_n30.t1 a_5452_n45.t5 VSS.t1973 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4042 a_3042_211.t1 RWLB[14].t12 a_2590_n953.t38 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4043 a_4192_3907.t0 VSS.t557 a_3740_n953.t10 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4044 a_3617_3425.t0 RWLB[1].t9 a_3165_n953.t31 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4045 VSS.t1518 a_4972_2421.t5 a_5342_2421.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4046 a_4767_1457.t1 RWLB[9].t14 a_4315_n953.t28 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4047 a_7177_4133.t2 WWLD[2].t26 a_7445_4887.t12 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4048 a_2672_211.t2 a_2577_196.t4 VDD.t1938 VDD.t1937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4049 a_2097_4686.t0 a_2002_4671.t5 VSS.t1811 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4050 a_3740_4445.t0 a_3727_4430.t5 VSS.t1055 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4051 a_6122_4445.t1 a_6027_4430.t5 VDD.t964 VDD.t963 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4052 a_5465_n953.t4 VSS.t556 a_5465_3907.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4053 a_8422_3907.t0 a_8327_3892.t4 VSS.t1447 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4054 a_6492_2943.t0 RWLB[3].t13 a_6040_n953.t35 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4055 VSS.t852 a_8997_2421.t5 a_8902_2406.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4056 a_3165_n953.t24 RWL[11].t10 a_3165_975.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4057 VDD.t466 a_4397_2180.t5 a_4302_2165.t1 VDD.t465 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4058 a_8997_1939.t1 a_8902_1924.t4 VSS.t925 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4059 VDD.t506 a_3247_4148.t5 a_3152_4133.t1 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4060 a_947_3907.t1 a_852_3892.t4 VSS.t888 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4061 a_6040_n30.t0 a_6027_n45.t5 VSS.t1751 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4062 a_14072_n4470.t0 VCLP.t92 a_13934_n4470.t1 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4063 a_2015_n953.t0 RWL[15].t13 a_2015_n30.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4064 VSS.t2123 a_7272_4148.t5 a_7642_4148.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4065 VSS.t885 a_8422_2180.t5 a_8792_2180.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4066 a_4408_n953.t15 WWL[4].t23 a_4397_2662.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4067 a_8327_2406.t2 WWL[5].t23 a_8595_4887.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4068 a_2015_n953.t11 VSS.t555 a_2015_n512.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4069 a_8327_n286.t1 WWLD[4].t22 a_8595_4887.t18 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4070 a_n52_n4483.t0 PRE_CLSA.t107 VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4071 VSS.t1242 a_2097_3907.t5 a_2002_3892.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4072 a_947_975.t2 a_852_960.t5 VSS.t850 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4073 a_4448_n5293.t1 VCLP.t93 a_4413_n5092.t0 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4074 a_2683_n953.t15 WWLD[2].t27 a_2672_4148.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4075 VDD.t1544 a_4972_1939.t5 a_4877_1924.t2 VDD.t1543 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4076 VSS.t1730 a_372_4148.t5 a_277_4133.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4077 a_4890_n953.t30 RWL[0].t15 a_4890_3666.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4078 a_7642_3907.t0 VSS.t554 a_7190_n953.t15 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4079 VDD.t798 a_2311_n5850.t3 ADC5_OUT[1].t1 VDD.t797 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4080 a_852_n1068.t0 WWLD[7].t24 a_1120_4887.t15 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4081 a_1427_3892.t0 WWLD[3].t25 a_1695_4887.t9 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4082 a_290_3425.t0 a_277_3410.t5 VSS.t2152 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4083 a_1440_3184.t0 a_1427_3169.t5 VSS.t861 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4084 a_1522_2662.t1 a_1427_2647.t5 VDD.t1409 VDD.t1408 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4085 VSS.t810 a_8997_1939.t4 a_9367_1939.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4086 a_5465_n953.t3 VSS.t553 a_5465_n271.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4087 a_5547_4686.t0 a_5452_4671.t4 VSS.t1405 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4088 a_8915_n953.t2 VSS.t552 a_8915_3907.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4089 a_4192_3425.t0 RWLB[1].t10 a_3740_n953.t3 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4090 a_3833_n953.t12 WWL[5].t24 a_3822_2421.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4091 a_6615_n953.t26 RWL[11].t11 a_6615_975.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4092 a_5630_n8026.t2 a_5857_n8583.t4 ADC8_OUT[3].t2 VSS.t1361 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4093 VSS.t780 a_5118_n2426.t0 a_5118_n2426.t1 VSS.t779 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4094 a_8902_n527.t0 WWLD[5].t27 a_9170_4887.t3 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4095 VSS.t1446 a_1522_3666.t5 a_1427_3651.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4096 a_5465_n953.t22 RWL[1].t13 a_5465_3425.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4097 a_8422_3425.t0 a_8327_3410.t4 VSS.t1417 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4098 a_6133_n953.t10 WWL[3].t23 a_6122_2943.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4099 a_8217_3666.t0 RWLB[0].t12 a_7765_n953.t29 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4100 a_9367_1698.t1 RWLB[8].t13 a_8915_n953.t46 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4101 a_4397_211.t2 a_4302_196.t4 VDD.t1534 VDD.t1533 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4102 a_947_3425.t1 a_852_3410.t4 VSS.t952 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4103 a_7994_n8026.t2 a_8221_n8583.t4 ADC10_OUT[3].t1 VSS.t243 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4104 a_3152_1683.t2 WWL[8].t25 a_3420_4887.t23 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4105 VSS.t2146 a_2097_n271.t5 a_2002_n286.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4106 a_7039_n8583.t2 ADC9_OUT[3].t4 VDD.t1980 VDD.t1979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4107 a_8340_4686.t1 a_8327_4671.t5 VSS.t1402 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4108 VSS.t1630 a_5547_3907.t5 a_5452_3892.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4109 a_3727_n1068.t0 WWLD[7].t25 a_3995_4887.t22 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4110 a_2672_n812.t2 a_2577_n827.t5 VDD.t984 VDD.t983 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4111 a_4302_678.t0 WWL[12].t24 a_4570_4887.t14 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4112 a_865_4686.t1 a_852_4671.t5 VSS.t1179 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4113 VSS.t1628 a_3247_975.t5 a_3152_960.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4114 VSS.t491 a_8997_211.t4 a_8902_196.t0 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4115 a_4972_4445.t2 a_4877_4430.t3 VSS.t2328 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4116 VSS.t821 a_2097_3425.t5 a_2002_3410.t2 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4117 VSS.t1197 a_6697_n1053.t4 a_6602_n1068.t1 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4118 a_4767_4686.t1 VSS.t551 a_4315_n953.t10 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4119 VDD.t490 a_8422_2421.t5 a_8327_2406.t1 VDD.t489 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4120 VSS.t948 a_3247_1698.t4 a_3617_1698.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4121 a_2097_2180.t2 a_2002_2165.t5 VDD.t914 VDD.t913 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 a_8915_n953.t8 VSS.t550 a_8915_n271.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4123 a_8792_1457.t1 RWLB[9].t15 a_8340_n953.t30 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4124 VDD.t1982 SA_OUT[12].t4 a_7210_n1371.t0 VDD.t1981 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4125 a_7642_3425.t0 RWLB[1].t11 a_7190_n953.t27 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 a_8291_n8071.t0 SAEN.t96 a_8488_n8026.t0 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4127 a_352_n2234.t1 Din[0].t1 VSS.t1244 VSS.t1243 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4128 a_1427_3410.t0 WWL[1].t26 a_1695_4887.t2 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4129 a_2577_1442.t0 WWL[9].t26 a_2845_4887.t13 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4130 VSS.t961 a_3247_n812.t4 a_3617_n812.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4131 a_7858_n953.t10 WWL[7].t26 a_7847_1939.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4132 a_8915_n953.t26 RWL[1].t14 a_8915_3425.t0 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4133 VDD.t1744 a_1522_3907.t5 a_1427_3892.t2 VDD.t1743 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4134 a_7190_n953.t24 RWL[11].t12 a_7190_975.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4135 a_2311_n7216.t0 PRE_CLSA.t108 VDD.t279 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4136 a_1440_n30.t0 a_1427_n45.t5 VSS.t1855 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4137 VSS.t1592 a_5547_n271.t5 a_5452_n286.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4138 VDD.t280 PRE_CLSA.t109 ADC5_OUT[1].t0 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4139 a_9367_1216.t1 RWLB[10].t13 a_8915_n953.t27 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4140 a_865_211.t1 a_852_196.t5 VSS.t1293 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4141 VDD.t367 a_7039_n4483.t4 ADC9_OUT[0].t2 VDD.t366 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4142 a_2672_3184.t2 a_2577_3169.t4 VSS.t2019 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4143 a_8433_n953.t21 WWL[4].t24 a_8422_2662.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4144 a_9405_n7216.t1 ADC11_OUT[2].t3 VDD.t2230 VDD.t1429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4145 VDD.t1073 SA_OUT[9].t4 a_5485_n1371.t2 VDD.t1072 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4146 a_6040_n953.t4 VSS.t549 a_6040_n512.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4147 a_3152_1201.t0 WWL[10].t26 a_3420_4887.t8 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4148 VDD.t2279 a_927_n2234.t4 a_1050_n2132.t1 VDD.t2278 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4149 VSS.t789 a_6122_3907.t5 a_6027_3892.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4150 VSS.t1869 a_6697_1457.t4 a_6602_1442.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4151 VSS.t1051 a_5547_3425.t5 a_5452_3410.t1 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4152 a_958_n953.t13 WWL[4].t25 a_947_2662.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4153 VSS.t44 a_3822_975.t5 a_3727_960.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4154 a_9367_211.t1 RWLB[14].t13 a_8915_n953.t40 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4155 a_4315_2662.t1 a_4302_2647.t4 VSS.t1228 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4156 VDD.t480 a_8997_1939.t5 a_8902_1924.t1 VDD.t479 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4157 a_290_n953.t31 RWL[8].t10 a_290_1698.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4158 a_1337_n7203.t0 VCLP.t94 a_1199_n7203.t1 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4159 VSS.t1606 a_2097_n512.t4 a_2467_n512.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4160 a_6027_678.t2 WWL[12].t25 a_6295_4887.t9 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4161 a_7283_n953.t6 WWL[12].t26 a_7272_693.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4162 VSS.t1312 a_3822_1698.t5 a_4192_1698.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4163 a_2590_4148.t1 a_2577_4133.t5 VSS.t1516 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4164 VSS.t2245 a_2672_3666.t5 a_3042_3666.t1 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4165 a_5547_2662.t1 a_5452_2647.t4 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4166 a_3727_1924.t0 WWL[7].t27 a_3995_4887.t18 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4167 VSS.t489 a_3247_1216.t4 a_3617_1216.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4168 a_4972_4148.t2 a_4877_4133.t4 VDD.t1687 VDD.t1686 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4169 a_9008_n953.t5 WWL[5].t25 a_8997_2421.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4170 a_3493_n4483.t0 PRE_CLSA.t110 VDD.t282 VDD.t281 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4171 a_290_n953.t11 VSS.t548 a_290_n812.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4172 a_7877_n1770.t0 SA_OUT[13].t4 a_7785_n1371.t2 VSS.t2033 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4173 VDD.t1525 a_1522_n271.t5 a_1427_n286.t2 VDD.t1524 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4174 a_11776_n7216.t2 ADC13_OUT[2].t4 a_11846_n7203.t0 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4175 VDD.t432 SA_OUT[14].t4 a_8360_n1371.t1 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4176 a_372_3184.t2 a_277_3169.t5 VDD.t644 VDD.t643 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4177 VDD.t498 a_3802_n2234.t4 a_3925_n2132.t1 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4178 VSS.t2179 a_3822_n812.t5 a_4192_n812.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4179 VDD.t1648 a_2672_975.t5 a_2577_960.t2 VDD.t1647 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4180 a_1892_3184.t0 RWLB[2].t13 a_1440_n953.t43 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4181 VSS.t2101 a_8568_n2426.t7 a_12701_n7825.t1 VSS.t2098 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4182 VDD.t1807 a_12963_n7216.t3 ADC14_OUT[2].t1 VDD.t565 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4183 a_5465_n812.t1 a_5452_n827.t5 VSS.t1961 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4184 VDD.t1689 a_1522_3425.t5 a_1427_3410.t2 VDD.t1688 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4185 a_2097_2662.t0 a_2002_2647.t5 VSS.t411 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4186 a_3740_2421.t0 a_3727_2406.t5 VSS.t914 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4187 a_6027_3651.t2 WWL[0].t24 a_6295_4887.t26 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4188 a_6122_2421.t1 a_6027_2406.t5 VDD.t670 VDD.t669 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4189 a_7177_1683.t0 WWL[8].t26 a_7445_4887.t0 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4190 a_5342_975.t0 RWLB[11].t15 a_4890_n953.t23 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4191 VSS.t1028 a_6122_n271.t5 a_6027_n286.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4192 a_n1460_n6503.t2 a_n1233_n7216.t4 ADC2_OUT[2].t2 VSS.t485 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4193 VSS.t2444 a_7847_n1053.t4 a_8217_n1053.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4194 a_2108_n953.t10 WWLD[3].t26 a_2097_3907.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4195 a_3740_n271.t1 a_3727_n286.t5 VSS.t1384 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4196 a_6122_n271.t1 a_6027_n286.t5 VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4197 a_n3792_n5293.t1 VCLP.t95 a_n3827_n5092.t0 VSS.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4198 a_5465_n953.t0 RWL[14].t14 a_5465_211.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4199 a_1695_4887.t6 PRE_SRAM.t38 VDD.t2077 VDD.t2076 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4200 VSS.t1873 a_7272_975.t5 a_7177_960.t1 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4201 VDD.t596 a_3247_1698.t5 a_3152_1683.t1 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4202 a_6615_452.t0 a_6602_437.t5 VSS.t1385 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4203 VDD.t1581 SA_OUT[11].t4 a_6635_n1371.t1 VDD.t1580 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4204 a_3258_n953.t23 WWLD[7].t26 a_3247_n1053.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4205 VSS.t1146 a_6122_3425.t5 a_6027_3410.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4206 VSS.t482 a_4397_211.t4 a_4302_196.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4207 VDD.t1532 a_2077_n2234.t4 a_2200_n2132.t1 VDD.t1531 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4208 VSS.t1150 a_5547_n512.t4 a_5917_n512.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4209 a_8792_4686.t0 VSS.t547 a_8340_n953.t6 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4210 VSS.t1149 a_7272_1698.t5 a_7642_1698.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4211 a_2577_4671.t0 WWLD[0].t26 a_2845_4887.t18 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4212 a_290_n953.t29 RWL[10].t12 a_290_1216.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4213 VDD.t604 a_3247_n812.t5 a_3152_n827.t2 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4214 a_8422_4148.t2 a_8327_4133.t5 VDD.t852 VDD.t851 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4215 a_7752_1442.t0 WWL[9].t27 a_8020_4887.t13 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4216 a_14072_n4470.t1 Iref0.t9 a_14131_n4114.t1 VSS.t2225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4217 a_1317_2180.t0 RWLB[6].t11 a_865_n953.t39 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4218 VDD.t1085 a_4675_n5850.t3 ADC7_OUT[1].t1 VDD.t1084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4219 a_1522_2943.t1 a_1427_2928.t5 VDD.t1234 VDD.t1233 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4220 VSS.t1721 a_3822_1216.t5 a_4192_1216.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4221 VSS.t1724 a_7272_n812.t5 a_7642_n812.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4222 a_1533_n953.t26 WWL[0].t25 a_1522_3666.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4223 a_2683_n953.t0 WWL[8].t27 a_2672_1698.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4224 VSS.t371 SAEN.t97 a_2084_n5293.t0 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4225 VSS.t1847 a_372_1698.t5 a_277_1683.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4226 VDD.t1298 a_4972_452.t5 a_4877_437.t2 VDD.t1297 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4227 a_9367_4445.t1 VSS.t546 a_8915_n953.t12 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4228 VSS.t2482 a_372_693.t5 a_277_678.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4229 VSS.t1154 a_6268_n2426.t0 a_6268_n2426.t1 VSS.t1153 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4230 a_8915_n812.t1 a_8902_n827.t4 VSS.t2198 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4231 a_5547_2662.t0 a_5452_2647.t5 VSS.t78 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4232 VSS.t2460 a_7847_1457.t4 a_8217_1457.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4233 a_7190_n953.t38 RWL[13].t12 a_7190_452.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4234 a_2108_n953.t13 WWLD[4].t23 a_2097_n271.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4235 a_18_n5338.t0 SAEN.t98 a_215_n5293.t0 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4236 a_2683_n953.t10 WWLD[6].t27 a_2672_n812.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4237 a_3152_4430.t2 WWLD[1].t26 a_3420_4887.t25 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4238 VDD.t874 a_4952_n2234.t4 a_5075_n2132.t1 VDD.t873 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4239 VSS.t912 a_372_n812.t5 a_277_n827.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4240 VSS.t1239 a_6697_4686.t4 a_6602_4671.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4241 a_10362_n8026.t2 a_10589_n8583.t4 ADC12_OUT[3].t2 VSS.t1564 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4242 VSS.t2327 a_6122_452.t5 a_6027_437.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4243 VDD.t2132 a_6697_452.t5 a_6602_437.t2 VDD.t2131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4244 VSS.t2130 a_7418_n2426.t0 a_7418_n2426.t1 VSS.t2129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4245 a_3258_n953.t14 WWL[9].t28 a_3247_1457.t2 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4246 a_7177_1201.t0 WWL[10].t27 a_7445_4887.t3 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4247 a_1522_n512.t0 a_1427_n527.t5 VSS.t46 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4248 a_2108_n953.t0 WWL[1].t27 a_2097_3425.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4249 a_6708_n953.t24 WWLD[7].t27 a_6697_n1053.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4250 VDD.t1348 a_2097_n512.t5 a_2002_n527.t1 VDD.t1347 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4251 VSS.t1728 a_3247_4445.t4 a_3617_4445.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4252 VDD.t1819 a_6122_3666.t5 a_6027_3651.t1 VDD.t1818 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4253 a_8340_2662.t0 a_8327_2647.t5 VSS.t1919 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4254 VDD.t424 a_3247_1216.t5 a_3152_1201.t2 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4255 a_4767_211.t1 RWLB[14].t14 a_4315_n953.t36 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4256 a_n3565_n5850.t1 ADC0_OUT[1].t3 VDD.t788 VDD.t364 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4257 a_3247_693.t0 a_3152_678.t5 VSS.t773 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4258 VSS.t1889 a_6122_n512.t5 a_6492_n512.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4259 a_6697_975.t2 a_6602_960.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4260 a_1427_678.t0 WWL[12].t27 a_1695_4887.t10 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4261 a_2683_n953.t5 WWL[12].t28 a_2672_693.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4262 a_6697_n812.t2 a_6602_n827.t5 VSS.t1617 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4263 a_865_2662.t0 a_852_2647.t5 VSS.t868 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4264 a_4972_2421.t1 a_4877_2406.t4 VSS.t2367 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4265 VSS.t1887 a_7272_1216.t5 a_7642_1216.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4266 a_156_n7203.t1 Iref2.t12 a_215_n6847.t1 VSS.t829 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4267 a_9613_n5338.t1 Iref1.t13 a_9672_n5293.t1 VSS.t2232 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4268 a_2015_n953.t33 EN.t11 a_n314_n4378.t0 VSS.t1951 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4269 a_6602_n1068.t2 WWLD[7].t28 a_6870_4887.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4270 a_7765_n512.t1 a_7752_n527.t5 VSS.t1743 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4271 a_4767_2662.t1 RWLB[4].t14 a_4315_n953.t34 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4272 a_4972_n271.t0 a_4877_n286.t4 VSS.t2354 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4273 a_277_1924.t2 WWL[7].t28 a_545_4887.t10 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4274 a_7067_3184.t0 RWLB[2].t14 a_6615_n953.t46 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4275 a_4972_693.t1 a_4877_678.t4 VSS.t1622 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4276 VSS.t1116 a_1522_n30.t5 a_1427_n45.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4277 a_7765_n30.t1 a_7752_n45.t5 VSS.t1165 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4278 a_852_3169.t2 WWL[2].t24 a_1120_4887.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4279 a_2683_n953.t3 WWL[10].t28 a_2672_1216.t1 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4280 a_3165_n953.t44 RWL[6].t11 a_3165_2180.t1 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4281 a_6122_2180.t1 a_6027_2165.t5 VSS.t2339 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4282 VSS.t394 a_372_1216.t5 a_277_1201.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4283 VDD.t1691 a_6697_975.t5 a_6602_960.t0 VDD.t1690 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4284 a_12963_n4483.t2 ADC14_OUT[0].t4 VDD.t1442 VDD.t1441 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4285 VDD.t2203 a_7847_n1053.t5 a_7752_n1068.t2 VDD.t2202 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4286 a_2015_n953.t3 VSS.t545 a_2015_4148.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4287 a_947_n30.t2 a_852_n45.t4 VDD.t1469 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4288 a_742_693.t1 RWLB[12].t12 a_290_n953.t20 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4289 a_372_211.t2 a_277_196.t4 VDD.t1672 VDD.t1671 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4290 a_3235_n1770.t2 PRE_VLSA.t42 VSS.t136 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4291 VDD.t824 a_372_n1053.t5 a_277_n1068.t1 VDD.t823 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4292 a_6133_n953.t6 WWLD[3].t27 a_6122_3907.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4293 a_6708_n953.t12 WWL[9].t29 a_6697_1457.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4294 a_6492_452.t0 RWLB[13].t12 a_6040_n953.t20 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4295 VDD.t779 a_5547_n512.t5 a_5452_n527.t1 VDD.t778 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 VSS.t2078 a_947_3184.t4 a_1317_3184.t0 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4297 a_1337_n4470.t0 VCLP.t96 a_1199_n4470.t1 VSS.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4298 a_290_n953.t14 VSS.t544 a_290_4445.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4299 a_2015_3907.t1 a_2002_3892.t4 VSS.t2120 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4300 a_n2345_n7203.t0 SAEN.t99 a_n2148_n6847.t0 VSS.t364 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4301 a_7283_n953.t13 WWLD[7].t29 a_7272_n1053.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4302 a_7752_4671.t0 WWLD[0].t27 a_8020_4887.t18 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4303 a_3420_4887.t14 WE.t28 a_3468_n2086.t0 VSS.t2411 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 VSS.t1053 a_3822_4445.t5 a_4192_4445.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4305 a_12736_n6503.t1 a_5743_n6391# a_12701_n6849.t0 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4306 a_4315_2943.t1 a_4302_2928.t4 VSS.t979 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4307 a_3247_3907.t2 a_3152_3892.t4 VDD.t2269 VDD.t2268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4308 a_7765_n953.t18 RWL[3].t15 a_7765_2943.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4309 a_2590_n953.t26 RWL[7].t14 a_2590_1939.t0 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4310 a_3822_1457.t1 a_3727_1442.t5 VDD.t1886 VDD.t1885 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4311 a_3701_n7203.t0 VCLP.t97 a_3563_n7203.t2 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4312 a_11776_n4483.t2 ADC13_OUT[0].t4 a_11846_n4470.t1 VSS.t862 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4313 a_4983_n953.t12 WWLD[5].t28 a_4972_n512.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4314 a_5547_2943.t1 a_5452_2928.t4 VDD.t2118 VDD.t2117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4315 a_5342_2180.t1 RWLB[6].t12 a_4890_n953.t25 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4316 a_3165_n953.t38 EN.t12 a_2049_n4378.t3 VSS.t1952 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4317 a_6110_n1770.t1 PRE_VLSA.t43 VSS.t140 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4318 VSS.t1673 a_7847_4686.t4 a_8217_4686.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4319 VDD.t2008 a_7847_1457.t5 a_7752_1442.t2 VDD.t2007 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4320 a_6615_n953.t45 RWL[6].t12 a_6615_2180.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4321 a_6065_n7203.t0 a_5743_n6391# a_5927_n7203.t2 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4322 VDD.t69 a_8422_n30.t5 a_8327_n45.t0 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4323 a_2590_1698.t1 a_2577_1683.t5 VSS.t2106 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4324 VDD.t1440 a_372_1457.t5 a_277_1442.t2 VDD.t1439 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4325 a_6133_n953.t17 WWLD[4].t24 a_6122_n271.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4326 a_n1460_n3770.t2 a_n1233_n4483.t4 ADC2_OUT[0].t2 VSS.t1837 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4327 a_3258_n953.t19 WWLD[0].t28 a_3247_4686.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4328 a_7177_4430.t0 WWLD[1].t27 a_7445_4887.t17 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4329 a_1440_3666.t0 a_1427_3651.t5 VSS.t1270 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4330 a_4972_1698.t0 a_4877_1683.t4 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4331 a_2590_n953.t39 RWL[13].t13 a_2590_452.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4332 VSS.t1357 a_4397_2943.t5 a_4302_2928.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4333 VSS.t1624 a_4972_693.t5 a_5342_693.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4334 a_290_n953.t2 RWL[15].t14 a_290_n30.t0 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4335 VSS.t1365 a_2097_n30.t5 a_2002_n45.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4336 a_8221_n4483.t0 PRE_CLSA.t111 VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4337 a_6295_4887.t12 WE.t29 a_6343_n2086.t0 VSS.t2412 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4338 a_2097_2943.t1 a_2002_2928.t5 VSS.t2028 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4339 VSS.t373 SAEN.t100 a_3266_n8026.t0 VSS.t372 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4340 VSS.t1533 a_1522_452.t5 a_1427_437.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4341 a_8997_n512.t1 a_8902_n527.t4 VSS.t1689 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4342 VDD.t1481 a_3247_4445.t5 a_3152_4430.t1 VDD.t1480 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4343 a_6133_n953.t0 WWL[1].t28 a_6122_3425.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4344 a_7283_n953.t14 WWL[9].t30 a_7272_1457.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4345 a_6122_452.t1 a_6027_437.t4 VDD.t2136 VDD.t2135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4346 a_4385_n1770.t0 PRE_VLSA.t44 VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4347 VSS.t388 a_3247_2180.t5 a_3152_2165.t1 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4348 VDD.t2079 PRE_SRAM.t39 a_958_n953.t23 VDD.t2078 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4349 VSS.t442 a_7272_4445.t5 a_7642_4445.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4350 a_3165_1457.t0 a_3152_1442.t5 VSS.t2046 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4351 a_n3357_n4470.t1 Iref0.t10 a_n3298_n4114.t1 VSS.t2226 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4352 a_6697_3907.t1 a_6602_3892.t5 VDD.t504 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4353 a_2015_3425.t1 a_2002_3410.t4 VSS.t1354 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4354 a_3420_4887.t5 PRE_SRAM.t40 a_3258_n953.t20 VDD.t2080 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4355 a_7847_452.t2 a_7752_437.t5 VDD.t2205 VDD.t2204 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4356 a_4570_4887.t24 WE.t30 a_4618_n2086.t1 VSS.t2413 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4357 a_2683_n953.t18 WWLD[1].t28 a_2672_4445.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4358 a_3247_3425.t1 a_3152_3410.t4 VDD.t1287 VDD.t1286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4359 a_2002_960.t0 WWL[11].t26 a_2270_4887.t3 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4360 a_5857_n7216.t1 ADC8_OUT[2].t4 a_5927_n7203.t0 VSS.t800 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4361 VSS.t2167 a_372_4445.t5 a_277_4430.t0 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4362 a_8792_2662.t0 RWLB[4].t15 a_8340_n953.t4 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4363 a_2577_2647.t2 WWL[4].t26 a_2845_4887.t8 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4364 a_2002_4133.t2 WWLD[2].t28 a_2270_4887.t19 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4365 a_4877_3169.t0 WWL[2].t25 a_5145_4887.t22 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4366 VSS.t374 SAEN.t101 a_4448_n5293.t0 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4367 a_6708_n953.t20 WWLD[0].t29 a_6697_4686.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4368 a_6040_n953.t3 VSS.t543 a_6040_4148.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4369 a_3247_3907.t1 a_3152_3892.t5 VSS.t2500 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4370 a_7190_n953.t44 RWL[6].t13 a_7190_2180.t0 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4371 VSS.t1425 a_2672_1939.t4 a_2577_1924.t2 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4372 a_8422_1698.t2 a_8327_1683.t5 VDD.t660 VDD.t659 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4373 a_9367_n1053.t0 VSS.t542 a_8915_n953.t1 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4374 a_3802_n2234.t1 Din[6].t1 VDD.t1354 VDD.t1353 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4375 VDD.t1825 a_947_3184.t5 a_852_3169.t1 VDD.t1824 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4376 a_5547_2943.t0 a_5452_2928.t5 VSS.t2293 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4377 a_2590_1216.t0 a_2577_1201.t5 VSS.t882 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4378 a_2311_n5850.t1 ADC5_OUT[1].t3 VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4379 a_4972_1216.t2 a_4877_1201.t4 VDD.t2172 VDD.t2171 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4380 a_9367_2421.t0 RWLB[5].t14 a_8915_n953.t18 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4381 VSS.t385 a_2097_4148.t4 a_2467_4148.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4382 a_1892_452.t1 RWLB[13].t13 a_1440_n953.t21 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4383 a_7752_196.t2 WWL[14].t27 a_8020_4887.t17 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4384 VSS.t812 a_4972_3184.t5 a_5342_3184.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4385 a_3152_2406.t2 WWL[5].t26 a_3420_4887.t12 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4386 a_7858_n953.t17 WWL[15].t27 a_7847_n30.t1 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4387 a_9367_n271.t0 VSS.t541 a_8915_n953.t13 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4388 a_7445_4887.t6 WE.t31 a_7493_n2086.t0 VSS.t2414 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 VSS.t2303 a_6697_2662.t4 a_6602_2647.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4390 a_383_n953.t2 WWL[11].t27 a_372_975.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4391 VDD.t285 PRE_CLSA.t112 ADC3_OUT[2].t0 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4392 a_3822_4686.t2 a_3727_4671.t5 VDD.t584 VDD.t583 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4393 a_6040_3907.t1 a_6027_3892.t5 VSS.t1343 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4394 VSS.t426 a_3822_2180.t5 a_3727_2165.t0 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4395 a_6615_1457.t0 a_6602_1442.t4 VSS.t815 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4396 a_3152_n286.t2 WWLD[4].t25 a_3420_4887.t15 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4397 VSS.t1206 a_8997_3184.t5 a_8902_3169.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4398 a_n279_n8026.t1 VCLP.t98 a_n314_n7825.t0 VSS.t176 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4399 a_8340_2943.t1 a_8327_2928.t5 VSS.t1380 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4400 a_2672_3666.t2 a_2577_3651.t5 VSS.t2332 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4401 a_7847_1457.t0 a_7752_1442.t4 VDD.t938 VDD.t937 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4402 VSS.t2047 a_372_n30.t5 a_277_n45.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4403 a_8221_n8583.t1 ADC10_OUT[3].t4 a_8291_n8071.t1 VSS.t246 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4404 VDD.t1411 a_7847_4686.t5 a_7752_4671.t2 VDD.t1410 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4405 a_6697_3425.t1 a_6602_3410.t5 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4406 a_2467_3907.t0 VSS.t540 a_2015_n953.t8 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4407 a_865_2943.t1 a_852_2928.t5 VSS.t1285 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4408 VDD.t1772 a_3822_2943.t5 a_3727_2928.t2 VDD.t1771 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4409 VSS.t1858 a_3247_2421.t4 a_3617_2421.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4410 a_6677_n2234.t1 Din[11].t1 VDD.t626 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4411 VDD.t632 a_372_4686.t5 a_277_4671.t0 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4412 a_5452_4133.t2 WWLD[2].t29 a_5720_4887.t21 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4413 a_8327_3169.t2 WWL[2].t26 a_8595_4887.t24 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4414 a_6602_2165.t2 WWL[6].t27 a_6870_4887.t6 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4415 a_7272_n30.t1 a_7177_n45.t4 VDD.t775 VDD.t774 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4416 a_742_4148.t0 VSS.t539 a_290_n953.t7 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4417 a_4767_2943.t0 RWLB[3].t14 a_4315_n953.t31 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4418 VDD.t1829 a_2672_2180.t5 a_2577_2165.t2 VDD.t1828 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4419 a_3727_960.t2 WWL[11].t28 a_3995_4887.t4 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4420 VDD.t1256 a_4397_n30.t5 a_4302_n45.t1 VDD.t1255 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4421 a_10797_n5338.t1 Iref1.t14 a_10856_n5293.t1 VSS.t2233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4422 a_3822_1939.t0 a_3727_1924.t5 VSS.t1551 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4423 a_4397_1457.t0 a_4302_1442.t5 VSS.t942 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4424 a_7283_n953.t22 WWLD[0].t30 a_7272_4686.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4425 a_3247_3425.t2 a_3152_3410.t5 VSS.t1535 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4426 VSS.t2127 a_8422_2943.t5 a_8327_2928.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4427 a_8422_1216.t2 a_8327_1201.t5 VDD.t1872 VDD.t1871 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4428 a_1440_n953.t15 VSS.t538 a_1440_n1053.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4429 VSS.t936 a_5547_4148.t4 a_5917_4148.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4430 a_372_3666.t2 a_277_3651.t5 VDD.t1946 VDD.t1945 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4431 a_7272_975.t2 a_7177_960.t5 VSS.t2036 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4432 a_3493_n8583.t2 ADC6_OUT[3].t4 VDD.t1181 VDD.t1180 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4433 a_n2345_n4470.t0 SAEN.t102 a_n2148_n4114.t0 VSS.t268 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4434 a_4952_n2234.t1 Din[8].t1 VDD.t846 VDD.t845 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4435 a_3165_4686.t1 a_3152_4671.t5 VSS.t1408 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4436 a_1892_3666.t1 RWLB[0].t13 a_1440_n953.t26 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4437 a_9008_n953.t4 WWL[12].t29 a_8997_693.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4438 VSS.t2475 a_7272_2180.t5 a_7177_2165.t2 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4439 a_2015_n953.t29 RWL[8].t11 a_2015_1698.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4440 a_1522_452.t1 a_1427_437.t5 VDD.t331 VDD.t330 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4441 a_12736_n3770.t1 VCLP.t99 a_12701_n4116.t0 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4442 VDD.t2082 PRE_SRAM.t41 a_4983_n953.t6 VDD.t2081 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4443 VSS.t2459 a_2049_n4378.t7 a_2049_n7825.t1 VSS.t2456 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4444 a_3833_n953.t3 WWL[2].t27 a_3822_3184.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4445 a_3701_n4470.t0 VCLP.t100 a_3563_n4470.t1 VSS.t203 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4446 a_6040_3425.t1 a_6027_3410.t5 VSS.t2088 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4447 a_8997_1939.t0 a_8902_1924.t5 VDD.t357 VDD.t356 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4448 a_7190_1457.t0 a_7177_1442.t5 VSS.t508 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 a_11984_n4470.t1 Iref0.t11 a_12043_n4114.t1 VSS.t2227 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4450 a_2015_n953.t6 VSS.t537 a_2015_n812.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4451 a_5917_3907.t0 VSS.t536 a_5465_n953.t10 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4452 a_290_n953.t48 RWL[5].t13 a_290_2421.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4453 a_7445_4887.t22 PRE_SRAM.t42 a_7283_n953.t24 VDD.t2083 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4454 a_7752_2647.t0 WWL[4].t27 a_8020_4887.t8 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4455 a_6065_n4470.t0 VCLP.t101 a_5927_n4470.t1 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4456 a_2467_3425.t1 RWLB[1].t12 a_2015_n953.t26 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4457 VSS.t873 a_3822_2421.t5 a_4192_2421.t0 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4458 VSS.t1219 a_7847_1939.t5 a_7752_1924.t1 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4459 VDD.t287 PRE_CLSA.t113 ADC9_OUT[3].t0 VDD.t286 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4460 a_7827_n2234.t1 Din[13].t1 VDD.t1242 VDD.t1241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4461 a_2590_4445.t0 a_2577_4430.t5 VSS.t1112 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4462 a_3727_n527.t0 WWLD[5].t29 a_3995_4887.t14 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4463 a_4972_4445.t0 a_4877_4430.t4 VDD.t57 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4464 a_7272_3907.t2 a_7177_3892.t5 VSS.t2196 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4465 a_4408_n953.t13 WWL[3].t24 a_4397_2943.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4466 a_1440_n953.t19 RWL[9].t14 a_1440_1457.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4467 a_7847_1457.t2 a_7752_1442.t5 VSS.t1782 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4468 a_1337_n4470.t1 Iref0.t12 a_1396_n4114.t1 VSS.t2228 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4469 VDD.t317 a_2097_4148.t5 a_2002_4133.t0 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4470 VDD.t79 a_8422_3184.t5 a_8327_3169.t1 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4471 VSS.t1798 a_7847_2662.t4 a_8217_2662.t1 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4472 a_8997_n30.t2 a_8902_n45.t5 VDD.t2232 VDD.t2231 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4473 a_13171_n5338.t1 Iref1.t15 a_13230_n5293.t1 VSS.t2234 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4474 VDD.t1246 a_4972_n30.t5 a_4877_n45.t1 VDD.t1245 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4475 a_2084_n5293.t2 a_2311_n5850.t4 ADC5_OUT[1].t2 VSS.t458 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4476 a_6615_4686.t1 a_6602_4671.t4 VSS.t1358 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4477 VDD.t1445 a_3493_n4483.t4 ADC6_OUT[0].t2 VDD.t1444 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4478 a_8902_n827.t0 WWLD[6].t28 a_9170_4887.t9 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4479 VSS.t2464 a_6122_4148.t5 a_6492_4148.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4480 a_7177_2406.t0 WWL[5].t27 a_7445_4887.t5 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4481 a_3152_196.t1 WWL[14].t28 a_3420_4887.t18 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4482 a_3833_n953.t22 WWL[15].t28 a_3822_n30.t0 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4483 VSS.t375 SAEN.t103 a_n279_n5293.t0 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4484 a_3258_n953.t9 WWL[4].t28 a_3247_2662.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4485 a_8915_n953.t21 RWL[14].t15 a_8915_211.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4486 a_7847_4686.t1 a_7752_4671.t4 VDD.t492 VDD.t491 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4487 a_7177_n286.t0 WWLD[4].t26 a_7445_4887.t18 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4488 a_2015_n953.t27 RWL[10].t13 a_2015_1216.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4489 a_9475_n5338.t0 SAEN.t104 a_9672_n5293.t0 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4490 VDD.t1614 a_3247_2421.t5 a_3152_2406.t1 VDD.t1613 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4491 a_6697_211.t1 a_6602_196.t5 VSS.t1371 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4492 a_5857_n4483.t1 ADC8_OUT[0].t4 a_5927_n4470.t2 VSS.t1444 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4493 a_4890_n1053.t1 a_4877_n1068.t5 VSS.t2365 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4494 a_2702_n1770.t0 SA_OUT[4].t4 a_2610_n1371.t2 VSS.t1704 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4495 a_6492_3907.t0 VSS.t535 a_6040_n953.t7 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4496 a_3042_n30.t1 RWLB[15].t13 a_2590_n953.t30 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4497 a_5917_3425.t1 RWLB[1].t13 a_5465_n953.t30 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4498 VSS.t2373 a_7272_2421.t5 a_7642_2421.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4499 a_4397_4686.t0 a_4302_4671.t5 VSS.t1852 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4500 a_8792_2943.t0 RWLB[3].t15 a_8340_n953.t32 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4501 a_5465_693.t1 a_5452_678.t5 VSS.t2277 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4502 a_2672_n30.t0 a_2577_n45.t5 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4503 a_n2207_n5338.t0 VCLP.t102 a_n2345_n5338.t2 VSS.t201 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4504 a_8915_n953.t45 EN.t13 a_8993_n2422.t0 VSS.t1953 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4505 a_8422_4445.t2 a_8327_4430.t5 VDD.t1642 VDD.t1641 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4506 a_7765_n953.t7 VSS.t534 a_7765_3907.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4507 a_383_n953.t9 WWL[12].t30 a_372_693.t0 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4508 a_2577_2928.t0 WWL[3].t25 a_2845_4887.t7 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4509 a_2683_n953.t6 WWL[5].t28 a_2672_2421.t2 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4510 a_5465_n953.t25 RWL[11].t13 a_5465_975.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4511 VSS.t902 a_7847_452.t5 a_7752_437.t0 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4512 a_10589_n7216.t1 ADC12_OUT[2].t4 a_10659_n7203.t1 VSS.t1530 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4513 VDD.t582 a_5547_4148.t5 a_5452_4133.t1 VDD.t581 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4514 VSS.t1675 a_372_2421.t5 a_277_2406.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4515 VDD.t9 a_6697_2180.t5 a_6602_2165.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4516 a_7272_3425.t2 a_7177_3410.t5 VSS.t1647 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4517 a_4877_437.t0 WWL[13].t27 a_5145_4887.t21 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4518 a_7190_211.t1 a_7177_196.t5 VSS.t1547 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4519 a_9613_n7203.t1 Iref2.t13 a_9672_n6847.t1 VSS.t830 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4520 a_7067_3666.t0 RWLB[0].t14 a_6615_n953.t30 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4521 a_6708_n953.t13 WWL[4].t29 a_6697_2662.t2 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4522 a_2002_1683.t0 WWL[8].t28 a_2270_4887.t0 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4523 VDD.t61 a_11776_n7216.t4 ADC13_OUT[2].t1 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4524 VSS.t910 a_352_n2234.t4 a_475_n2132.t0 VSS.t909 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4525 VDD.t2110 SA_OUT[2].t4 a_1460_n1371.t1 VDD.t2109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4526 a_4315_n953.t8 VSS.t533 a_4315_n512.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4527 a_7190_4686.t1 a_7177_4671.t5 VSS.t1526 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4528 a_852_3651.t2 WWL[0].t26 a_1120_4887.t23 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4529 VDD.t1448 a_n2415_n8583.t4 ADC1_OUT[3].t1 VDD.t1447 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4530 VSS.t1470 a_4397_3907.t5 a_4302_3892.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4531 a_9008_n953.t25 WWL[2].t28 a_8997_3184.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4532 a_6040_n953.t33 RWL[8].t12 a_6040_1698.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4533 a_2672_975.t1 a_2577_960.t5 VSS.t1738 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4534 a_4408_n953.t7 WWL[12].t31 a_4397_693.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4535 VSS.t1177 a_2097_975.t5 a_2002_960.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4536 VSS.t377 SAEN.t105 a_13637_n8026.t0 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4537 VSS.t2296 a_1522_n1053.t5 a_1892_n1053.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4538 a_4983_n953.t15 WWLD[2].t30 a_4972_4148.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4539 VDD.t1800 a_7272_1939.t5 a_7177_1924.t2 VDD.t1799 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4540 a_1129_n8583.t0 PRE_CLSA.t114 VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4541 a_7039_n5850.t1 ADC9_OUT[1].t3 VDD.t1674 VDD.t1673 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4542 a_4408_n953.t16 WWL[15].t29 a_4397_n30.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4543 a_n1233_n7216.t1 ADC2_OUT[2].t4 VDD.t2277 VDD.t1775 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4544 a_6040_n953.t13 VSS.t532 a_6040_n812.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4545 a_8217_1939.t0 RWLB[7].t13 a_7765_n953.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4546 a_6133_n953.t18 WWL[14].t29 a_6122_211.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4547 VSS.t1387 a_947_3666.t4 a_1317_3666.t1 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4548 a_3740_3184.t1 a_3727_3169.t5 VSS.t2002 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4549 a_3822_2662.t1 a_3727_2647.t5 VDD.t954 VDD.t953 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4550 VSS.t2479 a_2097_1698.t4 a_2467_1698.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4551 a_9178_n8026.t2 a_9405_n8583.t4 ADC11_OUT[3].t2 VSS.t1440 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4552 a_6122_3184.t2 a_6027_3169.t5 VDD.t749 VDD.t748 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4553 a_947_2180.t0 a_852_2165.t4 VDD.t658 VDD.t657 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4554 VSS.t2056 a_3247_n30.t5 a_3617_n30.t1 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4555 a_7765_n953.t12 VSS.t531 a_7765_n271.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4556 VSS.t1337 a_947_n512.t5 a_852_n527.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4557 a_1440_n953.t9 VSS.t530 a_1440_4686.t0 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4558 a_7847_4686.t0 a_7752_4671.t5 VSS.t833 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4559 a_3852_n1770.t0 SA_OUT[6].t4 a_3760_n1371.t1 VSS.t1427 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4560 a_6492_3425.t1 RWLB[1].t14 a_6040_n953.t29 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4561 VSS.t469 a_372_1939.t5 a_742_1939.t0 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 a_8915_n953.t23 RWL[11].t14 a_8915_975.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4563 VSS.t430 a_6697_211.t5 a_7067_211.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4564 VDD.t1548 a_7847_2662.t5 a_7752_2647.t2 VDD.t1547 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4565 a_8422_211.t2 a_8327_196.t5 VSS.t1908 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4566 a_10589_n7216.t0 PRE_CLSA.t115 VDD.t290 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4567 VSS.t460 a_2097_n812.t4 a_2467_n812.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4568 a_8433_n953.t18 WWL[3].t26 a_8422_2943.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4569 a_7765_n953.t22 RWL[1].t15 a_7765_3425.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4570 a_8217_452.t0 RWLB[13].t14 a_7765_n953.t21 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4571 VDD.t1075 a_372_2662.t5 a_277_2647.t1 VDD.t1074 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4572 a_277_n527.t0 WWLD[5].t30 a_545_4887.t4 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4573 a_3740_n953.t34 EN.t14 a_3231_n4378.t2 VSS.t1954 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4574 a_958_n953.t11 WWL[3].t27 a_947_2943.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4575 a_4397_n30.t2 a_4302_n45.t5 VDD.t606 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4576 a_5452_1683.t0 WWL[8].t29 a_5720_4887.t0 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4577 a_742_1698.t1 RWLB[8].t14 a_290_n953.t28 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4578 VSS.t1264 a_8422_211.t5 a_8792_211.t0 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4579 VDD.t1350 a_947_n30.t5 a_852_n45.t2 VDD.t1349 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4580 VSS.t1134 a_4397_n271.t5 a_4302_n286.t0 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4581 a_2015_n953.t12 VSS.t529 a_2015_4445.t0 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4582 VSS.t1204 a_1522_1457.t5 a_1892_1457.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4583 a_n2415_n4483.t2 ADC1_OUT[0].t4 VDD.t1071 VDD.t1070 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4584 a_7283_n953.t15 WWL[4].t30 a_7272_2662.t2 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4585 VSS.t791 a_5547_975.t5 a_5452_960.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4586 a_2002_1201.t2 WWL[10].t29 a_2270_4887.t5 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4587 a_290_n953.t40 RWL[13].t14 a_290_452.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4588 VSS.t2053 a_4397_3425.t5 a_4302_3410.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4589 a_6040_n953.t30 RWL[10].t14 a_6040_1216.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4590 a_3165_2662.t1 a_3152_2647.t5 VSS.t1718 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4591 VSS.t500 a_5547_1698.t4 a_5917_1698.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4592 VSS.t161 a_n3827_n4378.t7 a_n3827_n4116.t1 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4593 a_4397_2180.t1 a_4302_2165.t5 VDD.t508 VDD.t507 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4594 VSS.t103 a_4393_n2422.t7 a_4413_n4116.t1 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4595 a_7752_2928.t0 WWL[3].t28 a_8020_4887.t7 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4596 VSS.t449 a_2097_1216.t4 a_2467_1216.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4597 VSS.t379 SAEN.t106 a_6812_n8026.t0 VSS.t378 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4598 VSS.t1633 a_5547_n812.t4 a_5917_n812.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4599 a_4315_n953.t37 RWL[13].t15 a_4315_452.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4600 VDD.t2221 a_3822_3907.t5 a_3727_3892.t2 VDD.t2220 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4601 VSS.t2051 a_3247_452.t5 a_3152_437.t0 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4602 VSS.t1937 a_5075_n2132.t2 a_5053_n2086.t0 VSS.t1936 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4603 VDD.t706 a_1522_975.t5 a_1427_960.t2 VDD.t705 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4604 a_2097_452.t1 a_2002_437.t5 VSS.t808 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4605 a_2590_211.t0 a_2577_196.t5 VSS.t1302 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4606 a_3701_n4470.t1 Iref0.t13 a_3760_n4114.t1 VSS.t2229 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4607 a_2590_2421.t0 a_2577_2406.t5 VSS.t932 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4608 a_865_n30.t1 a_852_n45.t5 VSS.t1716 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4609 a_4877_3651.t2 WWL[0].t27 a_5145_4887.t23 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4610 a_4972_3184.t0 a_4877_3169.t4 VSS.t440 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4611 a_4972_2421.t2 a_4877_2406.t5 VDD.t2170 VDD.t2169 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4612 a_5452_1201.t0 WWL[10].t30 a_5720_4887.t6 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4613 a_2590_n271.t1 a_2577_n286.t5 VSS.t1196 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4614 a_4890_n953.t42 EN.t15 a_5118_n2426.t2 VSS.t1955 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4615 VSS.t1198 a_6697_n1053.t5 a_7067_n1053.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4616 a_8340_n953.t18 VSS.t528 a_8340_n512.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4617 a_4972_n271.t1 a_4877_n286.t5 VDD.t2162 VDD.t2161 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4618 VDD.t1530 a_n52_n7216.t4 ADC3_OUT[2].t2 VDD.t877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4619 a_4448_n5293.t2 a_4675_n5850.t4 ADC7_OUT[1].t2 VSS.t1224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4620 VSS.t413 a_8422_3907.t5 a_8327_3892.t1 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4621 a_742_1216.t1 RWLB[10].t14 a_290_n953.t38 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4622 a_865_n953.t15 VSS.t527 a_865_n512.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4623 a_902_n6503.t1 a_1129_n7216.t4 ADC4_OUT[2].t1 VSS.t1045 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4624 a_383_n953.t5 WWL[6].t28 a_372_2180.t2 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4625 VDD.t2242 a_2097_1698.t5 a_2002_1683.t1 VDD.t2241 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4626 VSS.t2473 a_6122_975.t5 a_6027_960.t2 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4627 a_6065_n4470.t1 Iref0.t14 a_6124_n4114.t1 VSS.t2230 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4628 VDD.t1021 a_947_3666.t5 a_852_3651.t1 VDD.t1020 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4629 a_6615_2662.t0 a_6602_2647.t5 VSS.t2261 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4630 a_9367_n30.t1 RWLB[15].t14 a_8915_n953.t43 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4631 VDD.t291 PRE_CLSA.t116 ADC6_OUT[2].t0 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4632 a_13864_n8583.t2 ADC15_OUT[3].t4 VDD.t1338 VDD.t1337 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4633 VSS.t446 a_3350_n2132.t2 a_3328_n2086.t0 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4634 VSS.t1044 a_4397_n512.t4 a_4767_n512.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4635 a_1129_n4483.t2 ADC4_OUT[0].t4 VDD.t1382 VDD.t1381 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4636 a_1522_n812.t1 a_1427_n827.t5 VSS.t878 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4637 VSS.t451 a_4972_3666.t5 a_5342_3666.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4638 a_7847_2662.t0 a_7752_2647.t4 VDD.t1507 VDD.t1506 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4639 VSS.t884 a_6122_1698.t5 a_6492_1698.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4640 VSS.t1581 a_5547_1216.t4 a_5917_1216.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4641 a_1533_n953.t19 WWL[14].t30 a_1522_211.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4642 a_4890_4148.t1 a_4877_4133.t5 VSS.t1912 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4643 a_6027_1924.t0 WWL[7].t29 a_6295_4887.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4644 VDD.t1107 PRE_VLSA.t45 a_6060_n1371.t0 VDD.t1106 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4645 VDD.t400 a_2097_n812.t5 a_2002_n827.t2 VDD.t399 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4646 VSS.t1110 a_4972_n512.t5 a_4877_n527.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4647 a_7272_4148.t2 a_7177_4133.t5 VDD.t1878 VDD.t1877 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4648 a_4972_693.t2 a_4877_678.t5 VDD.t1362 VDD.t1361 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4649 a_2577_n1068.t2 WWLD[7].t30 a_2845_4887.t23 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4650 VSS.t1626 a_8997_3666.t5 a_8902_3651.t1 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4651 a_5452_960.t0 WWL[11].t29 a_5720_4887.t3 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4652 VDD.t1426 a_3822_n271.t5 a_3727_n286.t2 VDD.t1425 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4653 a_10659_n5338.t0 SAEN.t107 a_10856_n5293.t0 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4654 VSS.t2024 a_2097_211.t5 a_2467_211.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4655 a_10589_n4483.t1 ADC12_OUT[0].t4 a_10659_n4470.t2 VSS.t1542 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4656 VSS.t1580 a_6122_n812.t5 a_6492_n812.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4657 a_3822_211.t1 a_3727_196.t5 VSS.t1187 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4658 a_n1025_n7203.t0 VCLP.t103 a_n1163_n7203.t1 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4659 a_3617_452.t0 RWLB[13].t15 a_3165_n953.t19 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4660 a_156_n7203.t0 VCLP.t104 a_18_n7203.t1 VSS.t218 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4661 a_n3565_n5850.t2 ADC0_OUT[1].t4 a_n3495_n5338.t2 VSS.t1164 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4662 a_7765_n812.t1 a_7752_n827.t5 VSS.t1140 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4663 VSS.t1636 a_1522_4686.t5 a_1892_4686.t1 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4664 VDD.t2267 a_3822_3425.t5 a_3727_3410.t2 VDD.t2266 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4665 a_4397_2662.t0 a_4302_2647.t5 VSS.t1229 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4666 a_8997_975.t0 a_8902_960.t5 VSS.t487 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4667 a_2002_4430.t2 WWLD[1].t29 a_2270_4887.t20 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4668 a_8422_2421.t1 a_8327_2406.t5 VDD.t888 VDD.t887 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4669 VSS.t1865 a_6697_1457.t5 a_7067_1457.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4670 a_4408_n953.t6 WWLD[3].t28 a_4397_3907.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4671 a_8327_3651.t2 WWL[0].t28 a_8595_4887.t15 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4672 VSS.t2010 a_8422_n271.t5 a_8327_n286.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4673 VDD.t293 PRE_CLSA.t117 ADC7_OUT[0].t0 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4674 VSS.t1700 a_6225_n2132.t2 a_6203_n2086.t1 VSS.t1699 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4675 a_6040_n953.t6 VSS.t526 a_6040_4445.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4676 a_2108_n953.t2 WWL[11].t30 a_2097_975.t2 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4677 a_8422_n271.t1 a_8327_n286.t5 VDD.t936 VDD.t935 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4678 VDD.t430 a_5547_1698.t5 a_5452_1683.t2 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4679 a_10797_n7203.t0 Iref2.t14 a_10856_n6847.t1 VSS.t831 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4680 a_6812_n5293.t1 VCLP.t105 a_6777_n5092.t0 VSS.t205 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4681 a_5558_n953.t19 WWLD[7].t31 a_5547_n1053.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4682 VSS.t1005 a_8422_3425.t5 a_8327_3410.t2 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4683 VDD.t862 a_13864_n4483.t4 ADC15_OUT[0].t2 VDD.t861 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4684 VSS.t1520 a_2097_4445.t4 a_2467_4445.t1 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4685 a_7190_2662.t0 a_7177_2647.t5 VSS.t1256 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4686 VDD.t389 a_2097_1216.t5 a_2002_1201.t0 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4687 VDD.t882 a_947_693.t5 a_852_678.t2 VDD.t881 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4688 VDD.t1376 a_5547_n812.t5 a_5452_n827.t2 VDD.t1375 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4689 a_1522_3907.t2 a_1427_3892.t5 VDD.t1865 VDD.t1864 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4690 VSS.t1452 a_3822_452.t5 a_4192_452.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4691 a_3822_2943.t2 a_3727_2928.t5 VDD.t1374 VDD.t1373 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4692 a_3617_2180.t0 RWLB[6].t13 a_3165_n953.t23 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4693 VSS.t765 a_6122_1216.t5 a_6492_1216.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4694 VSS.t1814 a_4500_n2132.t2 a_4478_n2086.t1 VSS.t1813 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4695 a_3833_n953.t26 WWL[0].t29 a_3822_3666.t2 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4696 a_4983_n953.t1 WWL[8].t30 a_4972_1698.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4697 VDD.t295 PRE_CLSA.t118 ADC2_OUT[0].t0 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4698 a_4192_n1053.t0 VSS.t525 a_3740_n953.t19 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4699 VDD.t1105 PRE_VLSA.t46 a_7210_n1371.t2 VDD.t1104 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4700 a_1440_n953.t45 RWL[4].t15 a_1440_2662.t1 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4701 a_7847_2662.t1 a_7752_2647.t5 VSS.t1767 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4702 a_4408_n953.t9 WWLD[4].t27 a_4397_n271.t2 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4703 a_13033_n5338.t0 SAEN.t108 a_13230_n5293.t0 VSS.t366 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4704 a_4983_n953.t0 WWLD[6].t29 a_4972_n812.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4705 a_5452_4430.t0 WWLD[1].t30 a_5720_4887.t22 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4706 VDD.t1455 a_5857_n7216.t4 ADC8_OUT[2].t2 VDD.t979 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4707 a_742_4445.t1 VSS.t524 a_290_n953.t8 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4708 a_4408_n953.t0 WWL[1].t29 a_4397_3425.t0 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4709 a_5558_n953.t20 WWL[9].t31 a_5547_1457.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4710 a_3822_n512.t0 a_3727_n527.t5 VSS.t57 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4711 a_6697_n1053.t0 a_6602_n1068.t5 VSS.t1910 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4712 VDD.t662 a_4397_n512.t5 a_4302_n527.t1 VDD.t661 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4713 VDD.t73 a_8221_n7216.t4 ADC10_OUT[2].t0 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4714 a_7272_n1053.t2 a_7177_n1068.t5 VDD.t1679 VDD.t1678 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4715 a_2467_n1053.t0 VSS.t523 a_2015_n953.t2 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4716 VSS.t1596 a_5547_4445.t4 a_5917_4445.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4717 VDD.t1415 a_8422_3666.t5 a_8327_3651.t1 VDD.t1414 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4718 VDD.t1328 a_5547_1216.t5 a_5452_1201.t2 VDD.t1327 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4719 a_2015_n953.t47 RWL[5].t14 a_2015_2421.t1 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4720 a_4767_n30.t1 RWLB[15].t15 a_4315_n953.t29 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4721 VSS.t970 a_8422_n512.t5 a_8792_n512.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4722 a_8997_n812.t0 a_8902_n827.t5 VSS.t2309 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4723 a_13171_n7203.t0 Iref2.t15 a_13230_n6847.t1 VSS.t832 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4724 a_3165_2943.t1 a_3152_2928.t5 VSS.t892 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4725 a_290_2180.t1 a_277_2165.t5 VSS.t484 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4726 a_1522_3425.t2 a_1427_3410.t5 VDD.t1837 VDD.t1836 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4727 a_2672_1457.t2 a_2577_1442.t5 VDD.t1732 VDD.t1731 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4728 a_n52_n8583.t2 ADC3_OUT[3].t4 a_18_n8071.t2 VSS.t1083 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4729 a_4675_n8583.t1 ADC7_OUT[3].t4 a_4745_n8071.t2 VSS.t1474 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4730 VSS.t496 a_3231_n4378.t7 a_3231_n5092.t1 VSS.t495 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4731 a_8997_n512.t2 a_8902_n527.t5 VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4732 a_3042_4148.t0 VSS.t522 a_2590_n953.t6 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4733 a_9367_3184.t1 RWLB[2].t15 a_8915_n953.t41 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4734 a_4192_2180.t0 RWLB[6].t14 a_3740_n953.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4735 a_4983_n953.t8 WWL[10].t31 a_4972_1216.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4736 a_6602_437.t0 WWL[13].t28 a_6870_4887.t18 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4737 VSS.t1240 a_6697_4686.t5 a_7067_4686.t1 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4738 a_3152_3169.t0 WWL[2].t29 a_3420_4887.t3 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4739 a_4315_n953.t7 VSS.t521 a_4315_4148.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4740 a_5465_n953.t45 RWL[6].t14 a_5465_2180.t1 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4741 a_8422_2180.t0 a_8327_2165.t5 VSS.t1060 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4742 a_13864_n8583.t0 PRE_CLSA.t119 VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4743 a_5342_n1053.t0 VSS.t520 a_4890_n953.t6 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4744 a_947_2180.t1 a_852_2165.t5 VSS.t1037 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4745 a_372_n30.t1 a_277_n45.t5 VDD.t678 VDD.t677 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4746 a_8433_n953.t10 WWLD[3].t29 a_8422_3907.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4747 VSS.t1928 a_n314_n4378.t7 a_n314_n5092.t1 VSS.t1922 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4748 a_902_n3770.t2 a_1129_n4483.t4 ADC4_OUT[0].t2 VSS.t1521 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4749 a_3165_975.t1 a_3152_960.t5 VSS.t1289 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4750 a_6133_n953.t23 WWL[11].t31 a_6122_975.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4751 a_958_n953.t5 WWLD[3].t30 a_947_3907.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4752 VSS.t1823 a_3247_3184.t4 a_3617_3184.t0 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4753 a_11984_n8071.t0 VCLP.t106 a_11846_n8071.t1 VSS.t224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4754 VDD.t1224 PRE_A.t15 a_5118_n2426.t3 VDD.t1223 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4755 VDD.t1269 a_2097_4445.t5 a_2002_4430.t1 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4756 a_7858_n953.t11 WWL[14].t31 a_7847_211.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4757 a_4315_3907.t1 a_4302_3892.t5 VSS.t1215 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4758 VSS.t1769 a_2097_2180.t5 a_2002_2165.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4759 a_n3792_n8026.t2 a_n3565_n8583.t4 ADC0_OUT[3].t2 VSS.t454 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4760 VSS.t1468 a_947_4148.t5 a_852_4133.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4761 VSS.t1252 a_6122_4445.t5 a_6492_4445.t1 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4762 a_6615_2943.t1 a_6602_2928.t5 VSS.t995 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4763 a_1440_1939.t0 a_1427_1924.t5 VSS.t1806 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4764 a_8422_n1053.t2 a_8327_n1068.t5 VDD.t698 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4765 a_7847_n1053.t1 a_7752_n1068.t5 VSS.t1161 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4766 a_5547_3907.t1 a_5452_3892.t4 VDD.t1585 VDD.t1584 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4767 a_4890_n953.t32 RWL[7].t15 a_4890_1939.t0 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4768 a_372_975.t2 a_277_960.t5 VSS.t1899 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4769 a_4890_975.t1 a_4877_960.t5 VSS.t2064 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4770 a_8291_n7203.t1 a_5632_n6430# a_8488_n6847.t0 VSS.t370 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4771 SA_OUT[8].t2 a_4910_n1371.t4 VDD.t1173 VDD.t1172 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4772 a_3617_n1053.t0 VSS.t519 a_3165_n953.t8 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4773 a_9008_n953.t17 WWL[0].t30 a_8997_3666.t2 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4774 a_n1460_n8026.t1 VCLP.t107 a_n1495_n7825.t0 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4775 a_2311_n5850.t2 ADC5_OUT[1].t4 a_2381_n5338.t2 VSS.t1126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4776 a_9405_n4483.t0 PRE_CLSA.t120 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4777 a_7642_2180.t0 RWLB[6].t15 a_7190_n953.t39 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4778 a_2270_4887.t25 PRE_SRAM.t43 a_2108_n953.t4 VDD.t2084 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4779 a_7847_2943.t2 a_7752_2928.t4 VDD.t1609 VDD.t1608 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4780 a_1427_2165.t0 WWL[6].t29 a_1695_4887.t11 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4781 a_n1025_n4470.t0 VCLP.t108 a_n1163_n4470.t1 VSS.t208 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4782 VDD.t300 PRE_CLSA.t121 ADC10_OUT[2].t2 VDD.t226 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4783 a_8915_n953.t36 RWL[6].t15 a_8915_2180.t1 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4784 a_8915_693.t1 a_8902_678.t5 VSS.t1121 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4785 a_156_n4470.t0 VCLP.t109 a_18_n4470.t1 VSS.t209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4786 a_2097_3907.t0 a_2002_3892.t5 VSS.t2121 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4787 a_3740_3666.t0 a_3727_3651.t5 VSS.t1185 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4788 a_4890_1698.t0 a_4877_1683.t5 VSS.t230 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4789 a_8433_n953.t13 WWLD[4].t28 a_8422_n271.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4790 a_5558_n953.t6 WWLD[0].t31 a_5547_4686.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4791 a_6122_3666.t1 a_6027_3651.t5 VDD.t1330 VDD.t1329 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4792 VSS.t804 a_6697_2943.t5 a_6602_2928.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4793 VSS.t837 a_1522_1939.t5 a_1427_1924.t1 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4794 a_7272_1698.t0 a_7177_1683.t5 VDD.t781 VDD.t780 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4795 a_2097_693.t1 a_2002_678.t5 VDD.t1652 VDD.t1651 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4796 a_958_n953.t19 WWLD[4].t29 a_947_n271.t2 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4797 SA_OUT[12].t2 a_7210_n1371.t4 a_7453_n1770.t0 VSS.t2048 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4798 SA_OUT[5].t2 a_3185_n1371.t4 VDD.t2195 VDD.t2194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4799 a_4397_2943.t1 a_4302_2928.t5 VSS.t980 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4800 a_8327_437.t0 WWL[13].t29 a_8595_4887.t23 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4801 VDD.t1344 a_5547_4445.t5 a_5452_4430.t2 VDD.t1343 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4802 a_372_4148.t1 a_277_4133.t5 VSS.t1319 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4803 a_290_n953.t0 RWL[2].t15 a_290_3184.t1 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4804 a_8433_n953.t0 WWL[1].t30 a_8422_3425.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4805 VSS.t1663 a_1522_2662.t5 a_1892_2662.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4806 VSS.t2006 a_3822_3184.t5 a_4192_3184.t1 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4807 VSS.t1330 a_5547_2180.t5 a_5452_2165.t2 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4808 VDD.t1428 a_7272_693.t5 a_7177_678.t1 VDD.t1427 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4809 a_7493_n2086.t1 a_7252_n2234.t4 VSS.t1503 VSS.t1502 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4810 a_958_n953.t0 WWL[1].t31 a_947_3425.t0 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4811 a_2002_2406.t0 WWL[5].t29 a_2270_4887.t8 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4812 VDD.t2086 PRE_SRAM.t44 a_3258_n953.t21 VDD.t2085 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4813 a_2672_4686.t1 a_2577_4671.t5 VDD.t1517 VDD.t1516 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4814 a_2002_n286.t0 WWLD[4].t30 a_2270_4887.t10 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4815 a_3810_n1770.t0 a_3995_4887.t27 a_4003_n1770.t0 VSS.t883 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4816 a_4315_3425.t1 a_4302_3410.t5 VSS.t1791 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4817 a_6040_n953.t47 RWL[5].t15 a_6040_2421.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4818 a_5465_1457.t0 a_5452_1442.t5 VSS.t1168 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4819 a_9405_n7216.t2 ADC11_OUT[2].t4 a_9475_n7203.t0 VSS.t2091 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4820 VDD.t1095 a_8997_211.t5 a_8902_196.t2 VDD.t1094 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4821 a_7190_2943.t1 a_7177_2928.t5 VSS.t1138 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4822 a_5720_4887.t26 PRE_SRAM.t45 a_5558_n953.t3 VDD.t2087 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4823 a_4983_n953.t23 WWLD[1].t31 a_4972_4445.t1 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4824 a_5547_3425.t1 a_5452_3410.t4 VDD.t1493 VDD.t1492 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4825 VSS.t492 a_8422_693.t5 a_8327_678.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4826 VDD.t301 PRE_CLSA.t122 ADC15_OUT[2].t0 VDD.t234 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4827 SA_OUT[9].t1 a_5485_n1371.t4 a_5728_n1770.t0 VSS.t498 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4828 VSS.t2145 a_2097_2421.t4 a_2467_2421.t0 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4829 a_7994_n6503.t1 a_5743_n6391# a_7959_n6849.t1 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4830 a_n2415_n8583.t0 PRE_CLSA.t123 VDD.t303 VDD.t302 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4831 SA_OUT[10].t1 a_6060_n1371.t4 VDD.t513 VDD.t512 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4832 a_8217_n512.t0 VSS.t518 a_7765_n953.t14 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4833 a_4302_4133.t1 WWLD[2].t31 a_4570_4887.t10 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4834 a_7177_3169.t0 WWL[2].t30 a_7445_4887.t25 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4835 a_5547_3907.t2 a_5452_3892.t5 VSS.t1833 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4836 a_8340_n953.t5 RWL[15].t15 a_8340_n30.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4837 a_8340_n953.t16 VSS.t517 a_8340_4148.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4838 VDD.t1384 a_1522_2180.t5 a_1427_2165.t1 VDD.t1383 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4839 a_2672_1939.t1 a_2577_1924.t5 VSS.t1835 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4840 a_865_n953.t16 VSS.t516 a_865_4148.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4841 a_2097_3425.t1 a_2002_3410.t5 VSS.t1355 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4842 VDD.t1575 a_3247_3184.t5 a_3152_3169.t2 VDD.t1574 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4843 a_7847_2943.t1 a_7752_2928.t5 VSS.t1854 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4844 a_4890_1216.t0 a_4877_1201.t5 VSS.t2368 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4845 a_6685_n1770.t0 a_6870_4887.t27 a_6878_n1770.t0 VSS.t1080 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4846 a_7272_1216.t0 a_7177_1201.t5 VDD.t554 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4847 a_4960_n1770.t2 PRE_VLSA.t47 VSS.t120 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4848 VSS.t2117 a_4397_4148.t4 a_4767_4148.t1 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4849 VSS.t1988 a_7272_3184.t5 a_7642_3184.t0 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4850 a_5452_2406.t0 WWL[5].t30 a_5720_4887.t9 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4851 a_7752_n45.t0 WWL[15].t30 a_8020_4887.t9 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4852 a_3727_n827.t0 WWLD[6].t30 a_3995_4887.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4853 VDD.t1509 a_10589_n7216.t4 ADC12_OUT[2].t2 VDD.t1508 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4854 a_12736_n6503.t2 a_12963_n7216.t4 ADC14_OUT[2].t2 VSS.t1538 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4855 SA_OUT[14].t2 a_8360_n1371.t4 a_8603_n1770.t0 VSS.t1481 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4856 SA_OUT[7].t2 a_4335_n1371.t4 VDD.t1177 VDD.t1176 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4857 a_8340_3907.t0 a_8327_3892.t5 VSS.t1448 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4858 a_742_2421.t0 RWLB[5].t15 a_290_n953.t47 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4859 a_8915_1457.t0 a_8902_1442.t5 VSS.t2165 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4860 a_7067_693.t0 RWLB[12].t13 a_6615_n953.t19 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4861 a_290_211.t1 a_277_196.t5 VSS.t1600 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4862 a_5452_n286.t2 WWLD[4].t31 a_5720_4887.t11 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4863 VSS.t1957 a_4972_4148.t5 a_4877_4133.t1 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4864 VSS.t1959 a_6122_2180.t5 a_6027_2165.t1 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4865 a_742_n271.t0 VSS.t515 a_290_n953.t4 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4866 VSS.t380 SAEN.t109 a_n1460_n5293.t0 VSS.t368 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4867 a_865_3907.t1 a_852_3892.t5 VSS.t889 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4868 a_4972_3666.t0 a_4877_3651.t5 VSS.t473 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4869 a_2683_n953.t25 WWL[2].t31 a_2672_3184.t0 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4870 a_3493_n5850.t2 ADC6_OUT[1].t4 VDD.t1192 VDD.t1054 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4871 a_8643_n2086.t0 a_8402_n2234.t4 VSS.t1011 VSS.t1010 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4872 VSS.t947 a_372_3184.t5 a_277_3169.t1 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4873 VDD.t1676 SA_OUT[0].t4 a_310_n1371.t2 VDD.t1675 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X4874 a_4767_3907.t0 VSS.t514 a_4315_n953.t9 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4875 a_6295_4887.t5 PRE_SRAM.t46 a_6133_n953.t22 VDD.t2088 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4876 VSS.t1336 a_5547_2421.t4 a_5917_2421.t1 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4877 a_372_1939.t1 a_277_1924.t5 VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4878 a_8792_693.t1 RWLB[12].t14 a_8340_n953.t23 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4879 VSS.t1254 a_7847_2943.t4 a_8217_2943.t0 VSS.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4880 VSS.t1426 a_2672_1939.t5 a_3042_1939.t0 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4881 a_1892_1939.t1 RWLB[7].t14 a_1440_n953.t0 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4882 a_4315_211.t1 a_4302_196.t5 VSS.t1786 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4883 a_3258_n953.t22 WWL[13].t30 a_3247_452.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4884 SA_OUT[11].t1 a_6635_n1371.t4 a_6878_n1770.t1 VSS.t921 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4885 a_3258_n953.t8 WWL[3].t29 a_3247_2943.t0 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4886 a_n3565_n8583.t0 PRE_CLSA.t124 VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4887 a_5547_3425.t2 a_5452_3410.t5 VSS.t1747 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4888 a_6697_1457.t0 a_6602_1442.t5 VSS.t816 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4889 VSS.t2096 a_8568_n2426.t0 a_8568_n2426.t1 VSS.t2095 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4890 a_3740_n953.t15 VSS.t513 a_3740_n1053.t0 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4891 VSS.t2300 a_6697_2662.t5 a_7067_2662.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4892 a_3042_1698.t1 RWLB[8].t15 a_2590_n953.t28 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4893 a_5547_452.t1 a_5452_437.t5 VSS.t1163 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4894 VDD.t306 PRE_CLSA.t125 ADC9_OUT[1].t0 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4895 a_3165_n953.t43 RWL[12].t14 a_3165_693.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4896 a_4983_n953.t18 WWL[13].t31 a_4972_452.t2 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4897 a_5465_4686.t0 a_5452_4671.t5 VSS.t1406 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4898 a_2108_n953.t5 WWL[6].t30 a_2097_2180.t0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4899 a_4315_n953.t30 RWL[8].t13 a_4315_1698.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4900 VSS.t944 a_2097_693.t5 a_2002_678.t1 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4901 VDD.t757 a_2672_693.t5 a_2577_678.t1 VDD.t756 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4902 VDD.t2090 PRE_SRAM.t47 a_7283_n953.t25 VDD.t2089 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4903 a_8291_n4470.t0 SAEN.t110 a_8488_n4114.t0 VSS.t279 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4904 a_8340_3425.t0 a_8327_3410.t5 VSS.t1752 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4905 a_9613_n7203.t0 a_5743_n6391# a_9475_n7203.t2 VSS.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4906 a_4315_n953.t3 VSS.t512 a_4315_n812.t0 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4907 VDD.t876 a_2097_2421.t5 a_2002_2406.t1 VDD.t875 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4908 a_4890_n953.t31 RWL[12].t15 a_4890_693.t1 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4909 a_6040_452.t0 a_6027_437.t5 VSS.t2263 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4910 VSS.t1508 a_3822_211.t5 a_3727_196.t2 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4911 VDD.t1029 a_4397_211.t5 a_4302_196.t2 VDD.t1028 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4912 a_865_3425.t1 a_852_3410.t5 VSS.t953 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4913 VSS.t1475 a_6122_2421.t5 a_6492_2421.t0 VSS.t260 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4914 a_4767_3425.t1 RWLB[1].t15 a_4315_n953.t26 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4915 VSS.t1594 a_947_1698.t5 a_852_1683.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4916 a_8422_693.t1 a_8327_678.t5 VDD.t538 VDD.t537 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4917 a_4890_4445.t1 a_4877_4430.t5 VSS.t2326 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4918 a_6708_n953.t11 WWL[3].t30 a_6697_2943.t0 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4919 a_1533_n953.t18 WWL[7].t30 a_1522_1939.t2 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4920 a_6027_n527.t2 WWLD[5].t31 a_6295_4887.t11 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4921 a_7272_4445.t2 a_7177_4430.t5 VDD.t1622 VDD.t1621 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4922 a_3740_n953.t22 RWL[9].t15 a_3740_1457.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4923 VSS.t107 a_5547_211.t5 a_5917_211.t0 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4924 VSS.t1400 a_8993_n2422.t7 a_13602_n5092.t1 VSS.t1394 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4925 a_7039_n5850.t2 ADC9_OUT[1].t4 a_7109_n5338.t2 VSS.t1504 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4926 VSS.t1758 a_947_n812.t5 a_852_n827.t2 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4927 VDD.t1870 a_4397_4148.t5 a_4302_4133.t2 VDD.t1869 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4928 a_8915_4686.t1 a_8902_4671.t5 VSS.t2522 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4929 VSS.t1900 a_8422_4148.t5 a_8792_4148.t1 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4930 a_3042_1216.t1 RWLB[10].t15 a_2590_n953.t37 VSS.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4931 a_5558_n953.t21 WWL[4].t31 a_5547_2662.t2 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4932 a_3152_n45.t0 WWL[15].t31 a_3420_4887.t22 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4933 a_3165_n953.t4 VSS.t511 a_3165_n512.t0 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4934 a_9405_n4483.t2 ADC11_OUT[0].t4 a_9475_n4470.t2 VSS.t905 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4935 a_2467_693.t0 RWLB[12].t15 a_2015_n953.t18 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4936 a_277_n827.t0 WWLD[6].t31 a_545_4887.t12 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4937 a_4315_n953.t0 RWL[10].t15 a_4315_1216.t1 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4938 a_8429_n8071.t0 VCLP.t110 a_8291_n8071.t2 VSS.t225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4939 VDD.t1839 a_5547_2421.t5 a_5452_2406.t2 VDD.t1838 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4940 VDD.t1813 a_6122_1939.t5 a_6027_1924.t2 VDD.t1812 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4941 a_156_n4470.t1 Iref0.t15 a_215_n4114.t1 VSS.t2231 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X4942 VDD.t880 a_7847_2943.t5 a_7752_2928.t2 VDD.t879 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4943 a_372_1698.t0 a_277_1683.t5 VSS.t1056 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4944 a_6697_n30.t2 a_6602_n45.t5 VSS.t1439 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4945 VDD.t1416 a_n2415_n5850.t4 ADC1_OUT[1].t2 VDD.t1044 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4946 a_7994_n3770.t1 VCLP.t111 a_7959_n4116.t0 VSS.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4947 a_8792_3907.t0 VSS.t510 a_8340_n953.t8 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4948 a_7067_1939.t0 RWLB[7].t15 a_6615_n953.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4949 a_4192_211.t0 RWLB[14].t15 a_3740_n953.t38 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4950 a_2577_3892.t0 WWLD[3].t31 a_2845_4887.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4951 a_2590_3184.t1 a_2577_3169.t5 VSS.t2020 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4952 VDD.t763 a_372_2943.t5 a_277_2928.t2 VDD.t762 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4953 a_2672_2662.t2 a_2577_2647.t5 VDD.t1587 VDD.t1586 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4954 a_852_1924.t2 WWL[7].t31 a_1120_4887.t10 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4955 VSS.t2197 a_7272_452.t5 a_7642_452.t1 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4956 a_4972_3184.t2 a_4877_3169.t5 VDD.t1754 VDD.t1753 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4957 a_1129_n5850.t0 PRE_CLSA.t126 VDD.t307 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4958 a_6697_4686.t0 a_6602_4671.t5 VSS.t1359 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4959 a_4983_n953.t11 WWL[5].t31 a_4972_2421.t0 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4960 VSS.t1836 a_947_1216.t5 a_852_1201.t1 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4961 a_7765_n953.t27 RWL[11].t15 a_7765_975.t0 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4962 a_7283_n953.t12 WWL[3].t31 a_7272_2943.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4963 VSS.t381 SAEN.t111 a_3266_n6503.t0 VSS.t372 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4964 a_7190_n30.t0 a_7177_n45.t5 VSS.t1929 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4965 a_12963_n4483.t0 PRE_CLSA.t127 VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X4966 a_9367_3666.t0 RWLB[0].t15 a_8915_n953.t30 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4967 a_12736_n3770.t2 a_12963_n4483.t4 ADC14_OUT[0].t1 VSS.t917 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=8e+06u l=150000u
X4968 a_3152_3651.t0 WWL[0].t31 a_3420_4887.t26 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4969 a_4302_1683.t0 WWL[8].t31 a_4570_4887.t2 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4970 a_6615_n953.t8 VSS.t509 a_6615_n512.t0 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4971 a_6133_n953.t2 WWL[6].t31 a_6122_2180.t0 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4972 VSS.t2297 a_6697_3907.t5 a_6602_3892.t0 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4973 a_8340_n953.t31 RWL[8].t14 a_8340_1698.t0 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4974 VSS.t2299 a_4397_975.t5 a_4302_960.t1 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4975 a_865_n953.t29 RWL[8].t15 a_865_1698.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 a_2002_2165.n0 a_2002_2165.t0 362.857
R1 a_2002_2165.t5 a_2002_2165.t4 337.399
R2 a_2002_2165.t4 a_2002_2165.t3 298.839
R3 a_2002_2165.n0 a_2002_2165.t5 280.405
R4 a_2002_2165.n1 a_2002_2165.t2 200
R5 a_2002_2165.n1 a_2002_2165.n0 172.311
R6 a_2002_2165.n2 a_2002_2165.n1 24
R7 a_2002_2165.n1 a_2002_2165.t1 21.212
R8 VSS.n339 VSS.t1947 3577.78
R9 VSS.n337 VSS.t1952 3511.11
R10 VSS.n342 VSS.t2043 3466.67
R11 VSS.n340 VSS.t1948 3422.22
R12 VSS.n336 VSS.t1951 3355.55
R13 VSS.n338 VSS.t1946 3355.55
R14 VSS.n335 VSS.t1945 3333.33
R15 VSS.n341 VSS.t1949 3311.11
R16 VSS.n341 VSS.t2042 3288.89
R17 VSS.n335 VSS.t1950 3266.67
R18 VSS.n336 VSS.t2044 3244.44
R19 VSS.n338 VSS.t1954 3244.44
R20 VSS.n340 VSS.t2041 3177.78
R21 VSS.n342 VSS.t1953 3133.33
R22 VSS.n337 VSS.t1944 3088.89
R23 VSS.n339 VSS.t1955 3022.22
R24 VSS.n2096 VSS.n2095 656.528
R25 VSS.n2092 VSS.n2091 637.705
R26 VSS.n2088 VSS.n2087 637.705
R27 VSS.n2084 VSS.n2083 637.705
R28 VSS.n2080 VSS.n2079 637.705
R29 VSS.n2076 VSS.n2075 637.705
R30 VSS.n2072 VSS.n2071 637.705
R31 VSS.n2068 VSS.n2067 637.705
R32 VSS.n2064 VSS.n2063 637.705
R33 VSS.n2060 VSS.n2059 637.705
R34 VSS.n2056 VSS.n2055 637.705
R35 VSS.n2052 VSS.n2051 637.705
R36 VSS.n2048 VSS.n2047 637.705
R37 VSS.n2044 VSS.n2043 637.705
R38 VSS.n2040 VSS.n2039 637.705
R39 VSS.n2036 VSS.n2035 637.705
R40 VSS.n2032 VSS.n2031 637.705
R41 VSS.n2290 VSS.t1366 616.124
R42 VSS.n2293 VSS.t1713 616.124
R43 VSS.n2296 VSS.t1485 616.124
R44 VSS.n2299 VSS.t1690 616.124
R45 VSS.n2302 VSS.t992 616.124
R46 VSS.n2305 VSS.t1368 616.124
R47 VSS.n2308 VSS.t2102 616.124
R48 VSS.n2311 VSS.t1222 616.124
R49 VSS.n2314 VSS.t2015 616.124
R50 VSS.n2317 VSS.t1614 616.124
R51 VSS.n2320 VSS.t1234 616.124
R52 VSS.n2323 VSS.t1282 616.124
R53 VSS.n2326 VSS.t1422 616.124
R54 VSS.n2329 VSS.t1759 616.124
R55 VSS.n2332 VSS.t2523 616.124
R56 VSS.n2290 VSS.t1008 560.113
R57 VSS.n2293 VSS.t402 560.113
R58 VSS.n2296 VSS.t1500 560.113
R59 VSS.n2299 VSS.t2066 560.113
R60 VSS.n2302 VSS.t865 560.113
R61 VSS.n2305 VSS.t1761 560.113
R62 VSS.n2308 VSS.t1245 560.113
R63 VSS.n2311 VSS.t1536 560.113
R64 VSS.n2314 VSS.t844 560.113
R65 VSS.n2317 VSS.t2506 560.113
R66 VSS.n2320 VSS.t1171 560.113
R67 VSS.n2323 VSS.t956 560.113
R68 VSS.n2326 VSS.t2274 560.113
R69 VSS.n2329 VSS.t2515 560.113
R70 VSS.n2332 VSS.t909 560.113
R71 VSS.n2289 VSS.t2401 498.131
R72 VSS.t2187 VSS.t2380 336.067
R73 VSS.t2192 VSS.t2392 336.067
R74 VSS.t76 VSS.t2379 336.067
R75 VSS.t2400 VSS.t2414 336.067
R76 VSS.t1080 VSS.t2393 336.067
R77 VSS.t1511 VSS.t2412 336.067
R78 VSS.t156 VSS.t2391 336.067
R79 VSS.t82 VSS.t2385 336.067
R80 VSS.t227 VSS.t2413 336.067
R81 VSS.t883 VSS.t2383 336.067
R82 VSS.t453 VSS.t2411 336.067
R83 VSS.t384 VSS.t2395 336.067
R84 VSS.t2423 VSS.t2384 336.067
R85 VSS.t1816 VSS.t2394 336.067
R86 VSS.t2267 VSS.t2382 336.067
R87 VSS.t2306 VSS.t2405 336.067
R88 VSS.n137 VSS.t278 327.137
R89 VSS.n128 VSS.t327 327.137
R90 VSS.n119 VSS.t369 327.137
R91 VSS.n110 VSS.t362 327.137
R92 VSS.n101 VSS.t317 327.137
R93 VSS.n92 VSS.t355 327.137
R94 VSS.n83 VSS.t265 327.137
R95 VSS.n74 VSS.t360 327.137
R96 VSS.n65 VSS.t307 327.137
R97 VSS.n56 VSS.t270 327.137
R98 VSS.n47 VSS.t310 327.137
R99 VSS.n38 VSS.t324 327.137
R100 VSS.n29 VSS.t314 327.137
R101 VSS.n20 VSS.t305 327.137
R102 VSS.n11 VSS.t295 327.137
R103 VSS.n2 VSS.t267 327.137
R104 VSS.n5 VSS.t283 327.137
R105 VSS.n14 VSS.t321 327.137
R106 VSS.n23 VSS.t328 327.137
R107 VSS.n32 VSS.t343 327.137
R108 VSS.n41 VSS.t349 327.137
R109 VSS.n50 VSS.t337 327.137
R110 VSS.n59 VSS.t288 327.137
R111 VSS.n68 VSS.t335 327.137
R112 VSS.n77 VSS.t374 327.137
R113 VSS.n86 VSS.t280 327.137
R114 VSS.n95 VSS.t371 327.137
R115 VSS.n104 VSS.t344 327.137
R116 VSS.n113 VSS.t375 327.137
R117 VSS.n122 VSS.t380 327.137
R118 VSS.n131 VSS.t353 327.137
R119 VSS.n331 VSS.t300 327.137
R120 VSS.n185 VSS.t263 327.137
R121 VSS.n182 VSS.t303 327.137
R122 VSS.n179 VSS.t351 327.137
R123 VSS.n176 VSS.t339 327.137
R124 VSS.n173 VSS.t293 327.137
R125 VSS.n170 VSS.t330 327.137
R126 VSS.n167 VSS.t373 327.137
R127 VSS.n164 VSS.t334 327.137
R128 VSS.n161 VSS.t285 327.137
R129 VSS.n158 VSS.t379 327.137
R130 VSS.n155 VSS.t287 327.137
R131 VSS.n152 VSS.t299 327.137
R132 VSS.n149 VSS.t290 327.137
R133 VSS.n146 VSS.t282 327.137
R134 VSS.n143 VSS.t274 327.137
R135 VSS.n140 VSS.t377 327.137
R136 VSS.n193 VSS.t1499 327.137
R137 VSS.n202 VSS.t1497 327.137
R138 VSS.n211 VSS.t1496 327.137
R139 VSS.n220 VSS.t1493 327.137
R140 VSS.n229 VSS.t1492 327.137
R141 VSS.n238 VSS.t1494 327.137
R142 VSS.n247 VSS.t1498 327.137
R143 VSS.n256 VSS.t1495 327.137
R144 VSS.n265 VSS.t356 327.137
R145 VSS.n274 VSS.t381 327.137
R146 VSS.n283 VSS.t352 327.137
R147 VSS.n292 VSS.t311 327.137
R148 VSS.n301 VSS.t358 327.137
R149 VSS.n310 VSS.t367 327.137
R150 VSS.n319 VSS.t319 327.137
R151 VSS.n328 VSS.t272 327.137
R152 VSS.t2164 VSS.t2404 317.397
R153 VSS.t2271 VSS.t2396 317.397
R154 VSS.t2301 VSS.t2390 317.397
R155 VSS.t2295 VSS.t2406 317.397
R156 VSS.t2305 VSS.t2389 317.397
R157 VSS.t6 VSS.t2403 317.397
R158 VSS.t968 VSS.t2410 317.397
R159 VSS.t2118 VSS.t2386 317.397
R160 VSS.t2304 VSS.t2398 317.397
R161 VSS.t455 VSS.t2388 317.397
R162 VSS.t2419 VSS.t2408 317.397
R163 VSS.t2166 VSS.t2399 317.397
R164 VSS.t2153 VSS.t2407 317.397
R165 VSS.t897 VSS.t2397 317.397
R166 VSS.t2178 VSS.t2387 317.397
R167 VSS.t2381 VSS.t803 317.397
R168 VSS.t1366 VSS.t2164 311.173
R169 VSS.t1713 VSS.t2271 311.173
R170 VSS.t1485 VSS.t2301 311.173
R171 VSS.t1690 VSS.t2295 311.173
R172 VSS.t992 VSS.t2305 311.173
R173 VSS.t1368 VSS.t6 311.173
R174 VSS.t2102 VSS.t968 311.173
R175 VSS.t1222 VSS.t2118 311.173
R176 VSS.t2015 VSS.t2304 311.173
R177 VSS.t1614 VSS.t455 311.173
R178 VSS.t1234 VSS.t2419 311.173
R179 VSS.t1282 VSS.t2166 311.173
R180 VSS.t1422 VSS.t2153 311.173
R181 VSS.t1759 VSS.t897 311.173
R182 VSS.t2523 VSS.t2178 311.173
R183 VSS.t133 VSS.t1902 311.173
R184 VSS.t803 VSS.t1243 311.173
R185 VSS.t2401 VSS.t2187 292.503
R186 VSS.t1008 VSS.t2192 292.503
R187 VSS.t402 VSS.t76 292.503
R188 VSS.t1500 VSS.t2400 292.503
R189 VSS.t2066 VSS.t1080 292.503
R190 VSS.t865 VSS.t1511 292.503
R191 VSS.t1761 VSS.t156 292.503
R192 VSS.t1245 VSS.t82 292.503
R193 VSS.t1536 VSS.t227 292.503
R194 VSS.t844 VSS.t883 292.503
R195 VSS.t2506 VSS.t453 292.503
R196 VSS.t1171 VSS.t384 292.503
R197 VSS.t956 VSS.t2423 292.503
R198 VSS.t2274 VSS.t1816 292.503
R199 VSS.t2515 VSS.t2267 292.503
R200 VSS.t909 VSS.t2306 292.503
R201 VSS.t2360 VSS.t143 280.056
R202 VSS.t1010 VSS.t129 280.056
R203 VSS.t405 VSS.t145 280.056
R204 VSS.t1502 VSS.t125 280.056
R205 VSS.t2068 VSS.t127 280.056
R206 VSS.t863 VSS.t139 280.056
R207 VSS.t1763 VSS.t123 280.056
R208 VSS.t1247 VSS.t119 280.056
R209 VSS.t972 VSS.t137 280.056
R210 VSS.t846 VSS.t121 280.056
R211 VSS.t2504 VSS.t135 280.056
R212 VSS.t1173 VSS.t147 280.056
R213 VSS.t1783 VSS.t141 280.056
R214 VSS.t801 VSS.t131 280.056
R215 VSS.t2512 VSS.t117 280.056
R216 VSS.t907 VSS.t133 280.056
R217 VSS.t2404 VSS.t2355 273.833
R218 VSS.t2396 VSS.t1280 273.833
R219 VSS.t2390 VSS.t395 273.833
R220 VSS.t2406 VSS.t1352 273.833
R221 VSS.t2389 VSS.t2115 273.833
R222 VSS.t2403 VSS.t1699 273.833
R223 VSS.t2410 VSS.t2017 273.833
R224 VSS.t2386 VSS.t1936 273.833
R225 VSS.t2398 VSS.t1813 273.833
R226 VSS.t2388 VSS.t949 273.833
R227 VSS.t2408 VSS.t445 273.833
R228 VSS.t2399 VSS.t1731 273.833
R229 VSS.t2407 VSS.t1642 273.833
R230 VSS.t2397 VSS.t1998 273.833
R231 VSS.t2387 VSS.t1693 273.833
R232 VSS.t937 VSS.t2381 273.833
R233 VSS.t2380 VSS.t978 261.386
R234 VSS.t2392 VSS.t1481 261.386
R235 VSS.t2379 VSS.t2034 261.386
R236 VSS.t2414 VSS.t2048 261.386
R237 VSS.t2393 VSS.t921 261.386
R238 VSS.t2412 VSS.t869 261.386
R239 VSS.t2391 VSS.t498 261.386
R240 VSS.t2385 VSS.t1458 261.386
R241 VSS.t2413 VSS.t1461 261.386
R242 VSS.t2383 VSS.t1565 261.386
R243 VSS.t2411 VSS.t2420 261.386
R244 VSS.t2395 VSS.t1122 261.386
R245 VSS.t2384 VSS.t399 261.386
R246 VSS.t2394 VSS.t154 261.386
R247 VSS.t2382 VSS.t1930 261.386
R248 VSS.t2405 VSS.t1464 261.386
R249 VSS.t181 VSS.t266 257.078
R250 VSS.t202 VSS.t294 257.078
R251 VSS.t183 VSS.t304 257.078
R252 VSS.t190 VSS.t313 257.078
R253 VSS.t171 VSS.t323 257.078
R254 VSS.t211 VSS.t309 257.078
R255 VSS.t205 VSS.t269 257.078
R256 VSS.t186 VSS.t306 257.078
R257 VSS.t192 VSS.t359 257.078
R258 VSS.t177 VSS.t264 257.078
R259 VSS.t189 VSS.t354 257.078
R260 VSS.t174 VSS.t316 257.078
R261 VSS.t179 VSS.t361 257.078
R262 VSS.t185 VSS.t368 257.078
R263 VSS.t180 VSS.t326 257.078
R264 VSS.t196 VSS.t277 257.078
R265 VSS.t200 VSS.t376 257.078
R266 VSS.t214 VSS.t273 257.078
R267 VSS.t206 VSS.t281 257.078
R268 VSS.t210 VSS.t289 257.078
R269 VSS.t223 VSS.t298 257.078
R270 VSS.t219 VSS.t286 257.078
R271 VSS.t178 VSS.t378 257.078
R272 VSS.t207 VSS.t284 257.078
R273 VSS.t164 VSS.t333 257.078
R274 VSS.t197 VSS.t372 257.078
R275 VSS.t163 VSS.t329 257.078
R276 VSS.t194 VSS.t292 257.078
R277 VSS.t176 VSS.t338 257.078
R278 VSS.t182 VSS.t350 257.078
R279 VSS.t199 VSS.t302 257.078
R280 VSS.t168 VSS.t262 257.078
R281 VSS.t59 VSS.t1236 239.775
R282 VSS.t1484 VSS.t917 239.775
R283 VSS.t862 VSS.t1856 239.775
R284 VSS.t1542 VSS.t1815 239.775
R285 VSS.t905 VSS.t1386 239.775
R286 VSS.t1698 VSS.t874 239.775
R287 VSS.t1504 VSS.t429 239.775
R288 VSS.t1444 VSS.t1341 239.775
R289 VSS.t1262 VSS.t1224 239.775
R290 VSS.t1181 VSS.t461 239.775
R291 VSS.t1126 VSS.t458 239.775
R292 VSS.t1638 VSS.t1521 239.775
R293 VSS.t900 VSS.t1837 239.775
R294 VSS.t494 VSS.t1676 239.775
R295 VSS.t1164 VSS.t427 239.775
R296 VSS.t1443 VSS.t1409 239.775
R297 VSS.t1540 VSS.t1538 239.775
R298 VSS.t87 VSS.t155 239.775
R299 VSS.t1530 VSS.t1564 239.775
R300 VSS.t2091 VSS.t1440 239.775
R301 VSS.t246 VSS.t243 239.775
R302 VSS.t1939 VSS.t991 239.775
R303 VSS.t800 VSS.t1361 239.775
R304 VSS.t1474 VSS.t1449 239.775
R305 VSS.t1424 VSS.t1376 239.775
R306 VSS.t1103 VSS.t1106 239.775
R307 VSS.t1046 VSS.t1045 239.775
R308 VSS.t1879 VSS.t485 239.775
R309 VSS.t1661 VSS.t1416 239.775
R310 VSS.t428 VSS.t454 239.775
R311 VSS.t195 VSS.t59 237.303
R312 VSS.t1236 VSS.t181 237.303
R313 VSS.t167 VSS.t1484 237.303
R314 VSS.t917 VSS.t202 237.303
R315 VSS.t184 VSS.t862 237.303
R316 VSS.t1856 VSS.t183 237.303
R317 VSS.t166 VSS.t1542 237.303
R318 VSS.t1815 VSS.t190 237.303
R319 VSS.t162 VSS.t905 237.303
R320 VSS.t1386 VSS.t171 237.303
R321 VSS.t187 VSS.t1698 237.303
R322 VSS.t874 VSS.t211 237.303
R323 VSS.t173 VSS.t1504 237.303
R324 VSS.t429 VSS.t205 237.303
R325 VSS.t204 VSS.t1444 237.303
R326 VSS.t1341 VSS.t186 237.303
R327 VSS.t172 VSS.t1262 237.303
R328 VSS.t1224 VSS.t192 237.303
R329 VSS.t203 VSS.t1181 237.303
R330 VSS.t461 VSS.t177 237.303
R331 VSS.t170 VSS.t1126 237.303
R332 VSS.t458 VSS.t189 237.303
R333 VSS.t198 VSS.t1638 237.303
R334 VSS.t1521 VSS.t174 237.303
R335 VSS.t209 VSS.t1123 237.303
R336 VSS.t1123 VSS.t1251 237.303
R337 VSS.t1251 VSS.t179 237.303
R338 VSS.t208 VSS.t900 237.303
R339 VSS.t1837 VSS.t185 237.303
R340 VSS.t201 VSS.t494 237.303
R341 VSS.t1676 VSS.t180 237.303
R342 VSS.t169 VSS.t1164 237.303
R343 VSS.t427 VSS.t196 237.303
R344 VSS.t212 VSS.t1443 237.303
R345 VSS.t1409 VSS.t200 237.303
R346 VSS.t222 VSS.t1540 237.303
R347 VSS.t1538 VSS.t214 237.303
R348 VSS.t224 VSS.t87 237.303
R349 VSS.t155 VSS.t206 237.303
R350 VSS.t221 VSS.t1530 237.303
R351 VSS.t1564 VSS.t210 237.303
R352 VSS.t220 VSS.t2091 237.303
R353 VSS.t1440 VSS.t223 237.303
R354 VSS.t225 VSS.t246 237.303
R355 VSS.t243 VSS.t219 237.303
R356 VSS.t193 VSS.t1939 237.303
R357 VSS.t991 VSS.t178 237.303
R358 VSS.t216 VSS.t800 237.303
R359 VSS.t1361 VSS.t207 237.303
R360 VSS.t191 VSS.t1474 237.303
R361 VSS.t1449 VSS.t164 237.303
R362 VSS.t215 VSS.t1424 237.303
R363 VSS.t1376 VSS.t197 237.303
R364 VSS.t188 VSS.t1103 237.303
R365 VSS.t1106 VSS.t163 237.303
R366 VSS.t213 VSS.t1046 237.303
R367 VSS.t1045 VSS.t194 237.303
R368 VSS.t218 VSS.t1083 237.303
R369 VSS.t1083 VSS.t96 237.303
R370 VSS.t96 VSS.t176 237.303
R371 VSS.t217 VSS.t1879 237.303
R372 VSS.t485 VSS.t182 237.303
R373 VSS.t175 VSS.t1661 237.303
R374 VSS.t1416 VSS.t199 237.303
R375 VSS.t165 VSS.t428 237.303
R376 VSS.t454 VSS.t168 237.303
R377 VSS.n0 VSS.t195 224.943
R378 VSS.n8 VSS.t167 224.943
R379 VSS.n17 VSS.t184 224.943
R380 VSS.n26 VSS.t166 224.943
R381 VSS.n35 VSS.t162 224.943
R382 VSS.n44 VSS.t187 224.943
R383 VSS.n53 VSS.t173 224.943
R384 VSS.n62 VSS.t204 224.943
R385 VSS.n71 VSS.t172 224.943
R386 VSS.n80 VSS.t203 224.943
R387 VSS.n89 VSS.t170 224.943
R388 VSS.n98 VSS.t198 224.943
R389 VSS.n107 VSS.t209 224.943
R390 VSS.n116 VSS.t208 222.471
R391 VSS.n125 VSS.t201 222.471
R392 VSS.n134 VSS.t169 222.471
R393 VSS.n6 VSS.n5 218.53
R394 VSS.n15 VSS.n14 218.53
R395 VSS.n24 VSS.n23 218.53
R396 VSS.n33 VSS.n32 218.53
R397 VSS.n42 VSS.n41 218.53
R398 VSS.n51 VSS.n50 218.53
R399 VSS.n60 VSS.n59 218.53
R400 VSS.n69 VSS.n68 218.53
R401 VSS.n78 VSS.n77 218.53
R402 VSS.n87 VSS.n86 218.53
R403 VSS.n96 VSS.n95 218.53
R404 VSS.n105 VSS.n104 218.53
R405 VSS.n114 VSS.n113 218.53
R406 VSS.n123 VSS.n122 218.53
R407 VSS.n132 VSS.n131 218.53
R408 VSS.n332 VSS.n331 218.53
R409 VSS.n186 VSS.n185 218.53
R410 VSS.n183 VSS.n182 218.53
R411 VSS.n180 VSS.n179 218.53
R412 VSS.n177 VSS.n176 218.53
R413 VSS.n174 VSS.n173 218.53
R414 VSS.n171 VSS.n170 218.53
R415 VSS.n168 VSS.n167 218.53
R416 VSS.n165 VSS.n164 218.53
R417 VSS.n162 VSS.n161 218.53
R418 VSS.n159 VSS.n158 218.53
R419 VSS.n156 VSS.n155 218.53
R420 VSS.n153 VSS.n152 218.53
R421 VSS.n150 VSS.n149 218.53
R422 VSS.n147 VSS.n146 218.53
R423 VSS.n144 VSS.n143 218.53
R424 VSS.n141 VSS.n140 218.53
R425 VSS.n194 VSS.n193 218.53
R426 VSS.n203 VSS.n202 218.53
R427 VSS.n212 VSS.n211 218.53
R428 VSS.n221 VSS.n220 218.53
R429 VSS.n230 VSS.n229 218.53
R430 VSS.n239 VSS.n238 218.53
R431 VSS.n248 VSS.n247 218.53
R432 VSS.n257 VSS.n256 218.53
R433 VSS.n266 VSS.n265 218.53
R434 VSS.n275 VSS.n274 218.53
R435 VSS.n284 VSS.n283 218.53
R436 VSS.n293 VSS.n292 218.53
R437 VSS.n302 VSS.n301 218.53
R438 VSS.n311 VSS.n310 218.53
R439 VSS.n320 VSS.n319 218.53
R440 VSS.n329 VSS.n328 218.53
R441 VSS.n189 VSS.t212 212.584
R442 VSS.n197 VSS.t222 212.584
R443 VSS.n206 VSS.t224 212.584
R444 VSS.n215 VSS.t221 212.584
R445 VSS.n224 VSS.t220 212.584
R446 VSS.n233 VSS.t225 212.584
R447 VSS.n242 VSS.t193 212.584
R448 VSS.n251 VSS.t216 212.584
R449 VSS.n260 VSS.t191 212.584
R450 VSS.n269 VSS.t215 212.584
R451 VSS.n278 VSS.t188 212.584
R452 VSS.n287 VSS.t213 212.584
R453 VSS.n296 VSS.t218 212.584
R454 VSS.n305 VSS.t217 210.112
R455 VSS.n314 VSS.t175 210.112
R456 VSS.n323 VSS.t165 210.112
R457 VSS.n2221 VSS.t1193 164.123
R458 VSS.n2218 VSS.t1963 164.123
R459 VSS.n2215 VSS.t2296 164.123
R460 VSS.n2212 VSS.t1378 164.123
R461 VSS.n2209 VSS.t2175 164.123
R462 VSS.n2206 VSS.t2169 164.123
R463 VSS.n2203 VSS.t2425 164.123
R464 VSS.n2200 VSS.t2442 164.123
R465 VSS.n2197 VSS.t2409 164.123
R466 VSS.n2194 VSS.t1996 164.123
R467 VSS.n2191 VSS.t1863 164.123
R468 VSS.n2188 VSS.t1198 164.123
R469 VSS.n2185 VSS.t1705 164.123
R470 VSS.n2182 VSS.t2444 164.123
R471 VSS.n2179 VSS.t1916 164.123
R472 VSS.n2177 VSS.t2193 164.123
R473 VSS.n1995 VSS.t2319 164.123
R474 VSS.n1992 VSS.t1225 164.123
R475 VSS.n1989 VSS.t1772 164.123
R476 VSS.n1986 VSS.t1606 164.123
R477 VSS.n1983 VSS.t2348 164.123
R478 VSS.n1980 VSS.t383 164.123
R479 VSS.n1977 VSS.t2362 164.123
R480 VSS.n1974 VSS.t1044 164.123
R481 VSS.n1971 VSS.t1109 164.123
R482 VSS.n1968 VSS.t1150 164.123
R483 VSS.n1965 VSS.t1889 164.123
R484 VSS.n1962 VSS.t2254 164.123
R485 VSS.n1959 VSS.t2160 164.123
R486 VSS.n1956 VSS.t1931 164.123
R487 VSS.n1953 VSS.t970 164.123
R488 VSS.n1951 VSS.t1740 164.123
R489 VSS.n1899 VSS.t2489 164.123
R490 VSS.n1896 VSS.t1567 164.123
R491 VSS.n1893 VSS.t1778 164.123
R492 VSS.n1890 VSS.t2151 164.123
R493 VSS.n1887 VSS.t1183 164.123
R494 VSS.n1884 VSS.t2199 164.123
R495 VSS.n1881 VSS.t1684 164.123
R496 VSS.n1878 VSS.t1880 164.123
R497 VSS.n1875 VSS.t971 164.123
R498 VSS.n1872 VSS.t1107 164.123
R499 VSS.n1869 VSS.t1027 164.123
R500 VSS.n1866 VSS.t77 164.123
R501 VSS.n1863 VSS.t2349 164.123
R502 VSS.n1860 VSS.t2249 164.123
R503 VSS.n1857 VSS.t2009 164.123
R504 VSS.n1855 VSS.t1098 164.123
R505 VSS.n1835 VSS.t1267 164.123
R506 VSS.n1832 VSS.t1607 164.123
R507 VSS.n1829 VSS.t1115 164.123
R508 VSS.n1826 VSS.t1364 164.123
R509 VSS.n1823 VSS.t239 164.123
R510 VSS.n1820 VSS.t2056 164.123
R511 VSS.n1817 VSS.t2209 164.123
R512 VSS.n1814 VSS.t1505 164.123
R513 VSS.n1811 VSS.t1488 164.123
R514 VSS.n1808 VSS.t1770 164.123
R515 VSS.n1805 VSS.t1709 164.123
R516 VSS.n1802 VSS.t1437 164.123
R517 VSS.n1799 VSS.t1843 164.123
R518 VSS.n1796 VSS.t1644 164.123
R519 VSS.n1793 VSS.t237 164.123
R520 VSS.n1791 VSS.t2477 164.123
R521 VSS.n1771 VSS.t1901 164.123
R522 VSS.n1768 VSS.t2241 164.123
R523 VSS.n1765 VSS.t1286 164.123
R524 VSS.n1762 VSS.t2024 164.123
R525 VSS.n1759 VSS.t1301 164.123
R526 VSS.n1756 VSS.t1599 164.123
R527 VSS.n1753 VSS.t1507 164.123
R528 VSS.n1750 VSS.t1801 164.123
R529 VSS.n1747 VSS.t1619 164.123
R530 VSS.n1744 VSS.t107 164.123
R531 VSS.n1741 VSS.t1260 164.123
R532 VSS.n1738 VSS.t430 164.123
R533 VSS.n1735 VSS.t152 164.123
R534 VSS.n1732 VSS.t1333 164.123
R535 VSS.n1729 VSS.t1264 164.123
R536 VSS.n1727 VSS.t490 164.123
R537 VSS.n1707 VSS.t2030 164.123
R538 VSS.n1704 VSS.t84 164.123
R539 VSS.n1701 VSS.t1660 164.123
R540 VSS.n1698 VSS.t1471 164.123
R541 VSS.n1695 VSS.t1529 164.123
R542 VSS.n1692 VSS.t1040 164.123
R543 VSS.n1689 VSS.t1452 164.123
R544 VSS.n1686 VSS.t437 164.123
R545 VSS.n1683 VSS.t1543 164.123
R546 VSS.n1680 VSS.t493 164.123
R547 VSS.n1677 VSS.t2324 164.123
R548 VSS.n1674 VSS.t2321 164.123
R549 VSS.n1671 VSS.t2197 164.123
R550 VSS.n1668 VSS.t448 164.123
R551 VSS.n1665 VSS.t1828 164.123
R552 VSS.n1663 VSS.t843 164.123
R553 VSS.n1562 VSS.t1588 164.123
R554 VSS.n1559 VSS.t797 164.123
R555 VSS.n1556 VSS.t996 164.123
R556 VSS.n1553 VSS.t1780 164.123
R557 VSS.n1550 VSS.t1883 164.123
R558 VSS.n1547 VSS.t1627 164.123
R559 VSS.n1544 VSS.t2376 164.123
R560 VSS.n1541 VSS.t2298 164.123
R561 VSS.n1538 VSS.t2000 164.123
R562 VSS.n1535 VSS.t772 164.123
R563 VSS.n1532 VSS.t2470 164.123
R564 VSS.n1529 VSS.t1915 164.123
R565 VSS.n1526 VSS.t1872 164.123
R566 VSS.n1523 VSS.t2514 164.123
R567 VSS.n1520 VSS.t2189 164.123
R568 VSS.n1518 VSS.t1268 164.123
R569 VSS.n1498 VSS.t401 164.123
R570 VSS.n1495 VSS.t1866 164.123
R571 VSS.n1492 VSS.t1552 164.123
R572 VSS.n1489 VSS.t449 164.123
R573 VSS.n1486 VSS.t1726 164.123
R574 VSS.n1483 VSS.t489 164.123
R575 VSS.n1480 VSS.t1721 164.123
R576 VSS.n1477 VSS.t2416 164.123
R577 VSS.n1474 VSS.t56 164.123
R578 VSS.n1471 VSS.t1581 164.123
R579 VSS.n1468 VSS.t765 164.123
R580 VSS.n1465 VSS.t1030 164.123
R581 VSS.n1462 VSS.t1887 164.123
R582 VSS.n1459 VSS.t792 164.123
R583 VSS.n1456 VSS.t2483 164.123
R584 VSS.n1454 VSS.t2060 164.123
R585 VSS.n1434 VSS.t1026 164.123
R586 VSS.n1431 VSS.t1189 164.123
R587 VSS.n1428 VSS.t1204 164.123
R588 VSS.n1425 VSS.t1679 164.123
R589 VSS.n1422 VSS.t1787 164.123
R590 VSS.n1419 VSS.t2073 164.123
R591 VSS.n1416 VSS.t875 164.123
R592 VSS.n1413 VSS.t1415 164.123
R593 VSS.n1410 VSS.t2216 164.123
R594 VSS.n1407 VSS.t1812 164.123
R595 VSS.n1404 VSS.t965 164.123
R596 VSS.n1401 VSS.t1865 164.123
R597 VSS.n1398 VSS.t1612 164.123
R598 VSS.n1395 VSS.t2460 164.123
R599 VSS.n1392 VSS.t1428 164.123
R600 VSS.n1390 VSS.t2302 164.123
R601 VSS.n1370 VSS.t1846 164.123
R602 VSS.n1367 VSS.t1593 164.123
R603 VSS.n1364 VSS.t1825 164.123
R604 VSS.n1361 VSS.t2479 164.123
R605 VSS.n1358 VSS.t1016 164.123
R606 VSS.n1355 VSS.t948 164.123
R607 VSS.n1352 VSS.t1312 164.123
R608 VSS.n1349 VSS.t389 164.123
R609 VSS.n1346 VSS.t1 164.123
R610 VSS.n1343 VSS.t500 164.123
R611 VSS.n1340 VSS.t884 164.123
R612 VSS.n1337 VSS.t1077 164.123
R613 VSS.n1334 VSS.t1149 164.123
R614 VSS.n1331 VSS.t1141 164.123
R615 VSS.n1328 VSS.t2168 164.123
R616 VSS.n1326 VSS.t2141 164.123
R617 VSS.n1306 VSS.t469 164.123
R618 VSS.n1303 VSS.t1061 164.123
R619 VSS.n1300 VSS.t836 164.123
R620 VSS.n1297 VSS.t2039 164.123
R621 VSS.n1294 VSS.t1426 164.123
R622 VSS.n1291 VSS.t1316 164.123
R623 VSS.n1288 VSS.t951 164.123
R624 VSS.n1285 VSS.t1857 164.123
R625 VSS.n1282 VSS.t1792 164.123
R626 VSS.n1279 VSS.t1682 164.123
R627 VSS.n1276 VSS.t1541 164.123
R628 VSS.n1273 VSS.t1809 164.123
R629 VSS.n1270 VSS.t2049 164.123
R630 VSS.n1267 VSS.t1218 164.123
R631 VSS.n1264 VSS.t1969 164.123
R632 VSS.n1262 VSS.t810 164.123
R633 VSS.n1242 VSS.t470 164.123
R634 VSS.n1239 VSS.t2143 164.123
R635 VSS.n1236 VSS.t1650 164.123
R636 VSS.n1233 VSS.t1768 164.123
R637 VSS.n1230 VSS.t2082 164.123
R638 VSS.n1227 VSS.t387 164.123
R639 VSS.n1224 VSS.t425 164.123
R640 VSS.n1221 VSS.t853 164.123
R641 VSS.n1218 VSS.t1942 164.123
R642 VSS.n1215 VSS.t1329 164.123
R643 VSS.n1212 VSS.t1958 164.123
R644 VSS.n1209 VSS.t49 164.123
R645 VSS.n1206 VSS.t2474 164.123
R646 VSS.n1203 VSS.t1669 164.123
R647 VSS.n1200 VSS.t885 164.123
R648 VSS.n1198 VSS.t2072 164.123
R649 VSS.n1178 VSS.t1674 164.123
R650 VSS.n1175 VSS.t2288 164.123
R651 VSS.n1172 VSS.t1681 164.123
R652 VSS.n1169 VSS.t2145 164.123
R653 VSS.n1166 VSS.t903 164.123
R654 VSS.n1163 VSS.t1858 164.123
R655 VSS.n1160 VSS.t873 164.123
R656 VSS.n1157 VSS.t1069 164.123
R657 VSS.n1154 VSS.t1518 164.123
R658 VSS.n1151 VSS.t1336 164.123
R659 VSS.n1148 VSS.t1475 164.123
R660 VSS.n1145 VSS.t1800 164.123
R661 VSS.n1142 VSS.t2373 164.123
R662 VSS.n1139 VSS.t890 164.123
R663 VSS.n1136 VSS.t822 164.123
R664 VSS.n1134 VSS.t851 164.123
R665 VSS.n1033 VSS.t1135 164.123
R666 VSS.n1030 VSS.t481 164.123
R667 VSS.n1027 VSS.t901 164.123
R668 VSS.n1024 VSS.t1232 164.123
R669 VSS.n1021 VSS.t2159 164.123
R670 VSS.n1018 VSS.t1002 164.123
R671 VSS.n1015 VSS.t2007 164.123
R672 VSS.n1012 VSS.t1356 164.123
R673 VSS.n1009 VSS.t927 164.123
R674 VSS.n1006 VSS.t835 164.123
R675 VSS.n1003 VSS.t1920 164.123
R676 VSS.n1000 VSS.t466 164.123
R677 VSS.n997 VSS.t1735 164.123
R678 VSS.n994 VSS.t1254 164.123
R679 VSS.n991 VSS.t2126 164.123
R680 VSS.n989 VSS.t1410 164.123
R681 VSS.n969 VSS.t1018 164.123
R682 VSS.n966 VSS.t2078 164.123
R683 VSS.n963 VSS.t1755 164.123
R684 VSS.n960 VSS.t2525 164.123
R685 VSS.n957 VSS.t2022 164.123
R686 VSS.n954 VSS.t1823 164.123
R687 VSS.n951 VSS.t2006 164.123
R688 VSS.n948 VSS.t1905 164.123
R689 VSS.n945 VSS.t812 164.123
R690 VSS.n942 VSS.t474 164.123
R691 VSS.n939 VSS.t1491 164.123
R692 VSS.n936 VSS.t1560 164.123
R693 VSS.n933 VSS.t1988 164.123
R694 VSS.n930 VSS.t1001 164.123
R695 VSS.n927 VSS.t234 164.123
R696 VSS.n925 VSS.t1205 164.123
R697 VSS.n905 VSS.t2272 164.123
R698 VSS.n902 VSS.t1803 164.123
R699 VSS.n899 VSS.t1913 164.123
R700 VSS.n896 VSS.t820 164.123
R701 VSS.n893 VSS.t1554 164.123
R702 VSS.n890 VSS.t2451 164.123
R703 VSS.n887 VSS.t2494 164.123
R704 VSS.n884 VSS.t2029 164.123
R705 VSS.n881 VSS.t1305 164.123
R706 VSS.n878 VSS.t1017 164.123
R707 VSS.n875 VSS.t1145 164.123
R708 VSS.n872 VSS.t2418 164.123
R709 VSS.n869 VSS.t478 164.123
R710 VSS.n866 VSS.t2204 164.123
R711 VSS.n863 VSS.t1004 164.123
R712 VSS.n861 VSS.t1088 164.123
R713 VSS.n841 VSS.t2207 164.123
R714 VSS.n838 VSS.t1387 164.123
R715 VSS.n835 VSS.t1445 164.123
R716 VSS.n832 VSS.t1989 164.123
R717 VSS.n829 VSS.t2245 164.123
R718 VSS.n826 VSS.t397 164.123
R719 VSS.n823 VSS.t40 164.123
R720 VSS.n820 VSS.t1586 164.123
R721 VSS.n817 VSS.t451 164.123
R722 VSS.n814 VSS.t1656 164.123
R723 VSS.n811 VSS.t2113 164.123
R724 VSS.n808 VSS.t1934 164.123
R725 VSS.n805 VSS.t2333 164.123
R726 VSS.n802 VSS.t1849 164.123
R727 VSS.n799 VSS.t465 164.123
R728 VSS.n797 VSS.t1625 164.123
R729 VSS.n745 VSS.t2320 164.123
R730 VSS.n742 VSS.t1390 164.123
R731 VSS.n739 VSS.t1788 164.123
R732 VSS.n736 VSS.t1241 164.123
R733 VSS.n733 VSS.t1891 164.123
R734 VSS.n730 VSS.t2370 164.123
R735 VSS.n727 VSS.t2446 164.123
R736 VSS.n724 VSS.t1469 164.123
R737 VSS.n721 VSS.t1748 164.123
R738 VSS.n718 VSS.t1629 164.123
R739 VSS.n715 VSS.t788 164.123
R740 VSS.n712 VSS.t2200 164.123
R741 VSS.n709 VSS.t2268 164.123
R742 VSS.n706 VSS.t2357 164.123
R743 VSS.n703 VSS.t412 164.123
R744 VSS.n701 VSS.t1867 164.123
R745 VSS.n574 VSS.t1729 164.123
R746 VSS.n577 VSS.t1467 164.123
R747 VSS.n580 VSS.t1413 164.123
R748 VSS.n583 VSS.t385 164.123
R749 VSS.n586 VSS.t1074 164.123
R750 VSS.n589 VSS.t859 164.123
R751 VSS.n592 VSS.t1081 164.123
R752 VSS.n595 VSS.t2117 164.123
R753 VSS.n598 VSS.t1956 164.123
R754 VSS.n601 VSS.t936 164.123
R755 VSS.n604 VSS.t2464 164.123
R756 VSS.n607 VSS.t2158 164.123
R757 VSS.n610 VSS.t2123 164.123
R758 VSS.n613 VSS.t1265 164.123
R759 VSS.n616 VSS.t1900 164.123
R760 VSS.n619 VSS.t2025 164.123
R761 VSS.n2094 VSS.t2208 164.123
R762 VSS.n1039 VSS.t906 164.123
R763 VSS.n1040 VSS.t1753 164.123
R764 VSS.n1043 VSS.t1663 164.123
R765 VSS.n1046 VSS.t1512 164.123
R766 VSS.n1049 VSS.t918 164.123
R767 VSS.n1052 VSS.t1372 164.123
R768 VSS.n1055 VSS.t1067 164.123
R769 VSS.n1058 VSS.t2031 164.123
R770 VSS.n1061 VSS.t2062 164.123
R771 VSS.n1064 VSS.t1124 164.123
R772 VSS.n1067 VSS.t1744 164.123
R773 VSS.n1070 VSS.t2300 164.123
R774 VSS.n1073 VSS.t418 164.123
R775 VSS.n1076 VSS.t1798 164.123
R776 VSS.n1079 VSS.t2075 164.123
R777 VSS.n1082 VSS.t1977 164.123
R778 VSS.n1566 VSS.t2481 164.123
R779 VSS.n1569 VSS.t1249 164.123
R780 VSS.n1572 VSS.t1294 164.123
R781 VSS.n1575 VSS.t943 164.123
R782 VSS.n1578 VSS.t1130 164.123
R783 VSS.n1581 VSS.t1831 164.123
R784 VSS.n1584 VSS.t251 164.123
R785 VSS.n1587 VSS.t2281 164.123
R786 VSS.n1590 VSS.t1624 164.123
R787 VSS.n1593 VSS.t149 164.123
R788 VSS.n1596 VSS.t1013 164.123
R789 VSS.n1599 VSS.t1087 164.123
R790 VSS.n1602 VSS.t1733 164.123
R791 VSS.n1605 VSS.t1658 164.123
R792 VSS.n1608 VSS.t1412 164.123
R793 VSS.n1611 VSS.t1118 164.123
R794 VSS.n2034 VSS.t911 164.123
R795 VSS.n2038 VSS.t1757 164.123
R796 VSS.n2042 VSS.t1462 164.123
R797 VSS.n2046 VSS.t460 164.123
R798 VSS.n2050 VSS.t1655 164.123
R799 VSS.n2054 VSS.t961 164.123
R800 VSS.n2058 VSS.t2179 164.123
R801 VSS.n2062 VSS.t158 164.123
R802 VSS.n2066 VSS.t111 164.123
R803 VSS.n2070 VSS.t1633 164.123
R804 VSS.n2074 VSS.t1580 164.123
R805 VSS.n2078 VSS.t1035 164.123
R806 VSS.n2082 VSS.t1724 164.123
R807 VSS.n2086 VSS.t2085 164.123
R808 VSS.n2090 VSS.t2215 164.123
R809 VSS.n536 VSS.t2337 164.123
R810 VSS.n533 VSS.t63 164.123
R811 VSS.n530 VSS.t1522 164.123
R812 VSS.n527 VSS.t1520 164.123
R813 VSS.n524 VSS.t946 164.123
R814 VSS.n521 VSS.t1728 164.123
R815 VSS.n518 VSS.t1053 164.123
R816 VSS.n515 VSS.t2428 164.123
R817 VSS.n512 VSS.t2426 164.123
R818 VSS.n509 VSS.t1596 164.123
R819 VSS.n506 VSS.t1252 164.123
R820 VSS.n503 VSS.t1712 164.123
R821 VSS.n500 VSS.t442 164.123
R822 VSS.n497 VSS.t1307 164.123
R823 VSS.n494 VSS.t1042 164.123
R824 VSS.n492 VSS.t1230 164.123
R825 VSS.n442 VSS.t1007 164.123
R826 VSS.n440 VSS.t1878 164.123
R827 VSS.n438 VSS.t1636 164.123
R828 VSS.n436 VSS.t839 164.123
R829 VSS.n434 VSS.t1777 164.123
R830 VSS.n432 VSS.t794 164.123
R831 VSS.n430 VSS.t1388 164.123
R832 VSS.n428 VSS.t1012 164.123
R833 VSS.n426 VSS.t2491 164.123
R834 VSS.n424 VSS.t414 164.123
R835 VSS.n422 VSS.t2111 164.123
R836 VSS.n420 VSS.t1240 164.123
R837 VSS.n418 VSS.t919 164.123
R838 VSS.n416 VSS.t1673 164.123
R839 VSS.n414 VSS.t1169 164.123
R840 VSS.n413 VSS.t2289 164.123
R841 VSS.n2272 VSS.t2466 162.724
R842 VSS.n2271 VSS.t964 162.724
R843 VSS.n2270 VSS.t1160 162.724
R844 VSS.n2269 VSS.t1904 162.724
R845 VSS.n2268 VSS.t1909 162.724
R846 VSS.n2267 VSS.t1876 162.724
R847 VSS.n2266 VSS.t767 162.724
R848 VSS.n2265 VSS.t2365 162.724
R849 VSS.n2264 VSS.t2445 162.724
R850 VSS.n2263 VSS.t2465 162.724
R851 VSS.n2262 VSS.t2186 162.724
R852 VSS.n2261 VSS.t2336 162.724
R853 VSS.n2260 VSS.t895 162.724
R854 VSS.n2259 VSS.t2308 162.724
R855 VSS.n2258 VSS.t1966 162.724
R856 VSS.n2257 VSS.t1192 162.724
R857 VSS.n2176 VSS.t2198 162.724
R858 VSS.n2175 VSS.t1460 162.724
R859 VSS.n2174 VSS.t1140 162.724
R860 VSS.n2173 VSS.t1720 162.724
R861 VSS.n2172 VSS.t1616 162.724
R862 VSS.n2171 VSS.t887 162.724
R863 VSS.n2170 VSS.t1961 162.724
R864 VSS.n2169 VSS.t226 162.724
R865 VSS.n2168 VSS.t2239 162.724
R866 VSS.n2167 VSS.t2247 162.724
R867 VSS.n2166 VSS.t959 162.724
R868 VSS.n2165 VSS.t1345 162.724
R869 VSS.n2164 VSS.t1310 162.724
R870 VSS.n2163 VSS.t877 162.724
R871 VSS.n2162 VSS.t1871 162.724
R872 VSS.n2161 VSS.t1079 162.724
R873 VSS.n1950 VSS.t1340 162.724
R874 VSS.n1949 VSS.t1297 162.724
R875 VSS.n1948 VSS.t2291 162.724
R876 VSS.n1947 VSS.t2352 162.724
R877 VSS.n1946 VSS.t113 162.724
R878 VSS.n1945 VSS.t1032 162.724
R879 VSS.n1944 VSS.t1144 162.724
R880 VSS.n1943 VSS.t2353 162.724
R881 VSS.n1942 VSS.t1084 162.724
R882 VSS.n1941 VSS.t1384 162.724
R883 VSS.n1940 VSS.t1877 162.724
R884 VSS.n1939 VSS.t1196 162.724
R885 VSS.n1938 VSS.t2149 162.724
R886 VSS.n1937 VSS.t2090 162.724
R887 VSS.n1936 VSS.t1570 162.724
R888 VSS.n1935 VSS.t2517 162.724
R889 VSS.n1854 VSS.t2476 162.724
R890 VSS.n1853 VSS.t247 162.724
R891 VSS.n1852 VSS.t1165 162.724
R892 VSS.n1851 VSS.t1929 162.724
R893 VSS.n1850 VSS.t1438 162.724
R894 VSS.n1849 VSS.t1751 162.724
R895 VSS.n1848 VSS.t1972 162.724
R896 VSS.n1847 VSS.t1490 162.724
R897 VSS.n1846 VSS.t423 162.724
R898 VSS.n1845 VSS.t2212 162.724
R899 VSS.n1844 VSS.t1971 162.724
R900 VSS.n1843 VSS.t110 162.724
R901 VSS.n1842 VSS.t1362 162.724
R902 VSS.n1841 VSS.t1855 162.724
R903 VSS.n1840 VSS.t1716 162.724
R904 VSS.n1839 VSS.t435 162.724
R905 VSS.n1790 VSS.t1058 162.724
R906 VSS.n1789 VSS.t1907 162.724
R907 VSS.n1788 VSS.t1332 162.724
R908 VSS.n1787 VSS.t1547 162.724
R909 VSS.n1786 VSS.t1370 162.724
R910 VSS.n1785 VSS.t1152 162.724
R911 VSS.n1784 VSS.t160 162.724
R912 VSS.n1783 VSS.t506 162.724
R913 VSS.n1782 VSS.t1786 162.724
R914 VSS.n1781 VSS.t1186 162.724
R915 VSS.n1780 VSS.t939 162.724
R916 VSS.n1779 VSS.t1302 162.724
R917 VSS.n1778 VSS.t1257 162.724
R918 VSS.n1777 VSS.t1895 162.724
R919 VSS.n1776 VSS.t1293 162.724
R920 VSS.n1775 VSS.t1600 162.724
R921 VSS.n1726 VSS.t841 162.724
R922 VSS.n1725 VSS.t923 162.724
R923 VSS.n1724 VSS.t2258 162.724
R924 VSS.n1723 VSS.t1108 162.724
R925 VSS.n1722 VSS.t1385 162.724
R926 VSS.n1721 VSS.t2263 162.724
R927 VSS.n1720 VSS.t1162 162.724
R928 VSS.n1719 VSS.t814 162.724
R929 VSS.n1718 VSS.t1314 162.724
R930 VSS.n1717 VSS.t1454 162.724
R931 VSS.n1716 VSS.t2054 162.724
R932 VSS.n1715 VSS.t1974 162.724
R933 VSS.n1714 VSS.t807 162.724
R934 VSS.n1713 VSS.t393 162.724
R935 VSS.n1712 VSS.t2431 162.724
R936 VSS.n1711 VSS.t443 162.724
R937 VSS.n1662 VSS.t1121 162.724
R938 VSS.n1661 VSS.t893 162.724
R939 VSS.n1660 VSS.t1327 162.724
R940 VSS.n1659 VSS.t2344 162.724
R941 VSS.n1658 VSS.t1099 162.724
R942 VSS.n1657 VSS.t975 162.724
R943 VSS.n1656 VSS.t2277 162.724
R944 VSS.n1655 VSS.t1621 162.724
R945 VSS.n1654 VSS.t2290 162.724
R946 VSS.n1653 VSS.t248 162.724
R947 VSS.n1652 VSS.t790 162.724
R948 VSS.n1651 VSS.t2499 162.724
R949 VSS.n1650 VSS.t1884 162.724
R950 VSS.n1649 VSS.t422 162.724
R951 VSS.n1648 VSS.t2469 162.724
R952 VSS.n1647 VSS.t2259 162.724
R953 VSS.n1517 VSS.t2014 162.724
R954 VSS.n1516 VSS.t504 162.724
R955 VSS.n1515 VSS.t787 162.724
R956 VSS.n1514 VSS.t1597 162.724
R957 VSS.n1513 VSS.t1774 162.724
R958 VSS.n1512 VSS.t1610 162.724
R959 VSS.n1511 VSS.t1562 162.724
R960 VSS.n1510 VSS.t2368 162.724
R961 VSS.n1509 VSS.t105 162.724
R962 VSS.n1508 VSS.t1664 162.724
R963 VSS.n1507 VSS.t998 162.724
R964 VSS.n1506 VSS.t882 162.724
R965 VSS.n1505 VSS.t799 162.724
R966 VSS.n1504 VSS.t1532 162.724
R967 VSS.n1503 VSS.t1478 162.724
R968 VSS.n1502 VSS.t390 162.724
R969 VSS.n1453 VSS.t2165 162.724
R970 VSS.n1452 VSS.t1114 162.724
R971 VSS.n1451 VSS.t1300 162.724
R972 VSS.n1450 VSS.t508 162.724
R973 VSS.n1449 VSS.t815 162.724
R974 VSS.n1448 VSS.t1583 162.724
R975 VSS.n1447 VSS.t1168 162.724
R976 VSS.n1446 VSS.t2210 162.724
R977 VSS.n1445 VSS.t941 162.724
R978 VSS.n1444 VSS.t2137 162.724
R979 VSS.n1443 VSS.t2046 162.724
R980 VSS.n1442 VSS.t1299 162.724
R981 VSS.n1441 VSS.t954 162.724
R982 VSS.n1440 VSS.t1202 162.724
R983 VSS.n1439 VSS.t2080 162.724
R984 VSS.n1438 VSS.t915 162.724
R985 VSS.n1389 VSS.t416 162.724
R986 VSS.n1388 VSS.t1039 162.724
R987 VSS.n1387 VSS.t2093 162.724
R988 VSS.n1386 VSS.t2140 162.724
R989 VSS.n1385 VSS.t1935 162.724
R990 VSS.n1384 VSS.t2125 162.724
R991 VSS.n1383 VSS.t1483 162.724
R992 VSS.n1382 VSS.t230 162.724
R993 VSS.n1381 VSS.t2252 162.724
R994 VSS.n1380 VSS.t1985 162.724
R995 VSS.n1379 VSS.t1652 162.724
R996 VSS.n1378 VSS.t2106 162.724
R997 VSS.n1377 VSS.t2467 162.724
R998 VSS.n1376 VSS.t1309 162.724
R999 VSS.n1375 VSS.t1591 162.724
R1000 VSS.n1374 VSS.t1668 162.724
R1001 VSS.n1325 VSS.t1473 162.724
R1002 VSS.n1324 VSS.t2237 162.724
R1003 VSS.n1323 VSS.t1807 162.724
R1004 VSS.n1322 VSS.t1701 162.724
R1005 VSS.n1321 VSS.t1381 162.724
R1006 VSS.n1320 VSS.t977 162.724
R1007 VSS.n1319 VSS.t1176 162.724
R1008 VSS.n1318 VSS.t58 162.724
R1009 VSS.n1317 VSS.t819 162.724
R1010 VSS.n1316 VSS.t1550 162.724
R1011 VSS.n1315 VSS.t1313 162.724
R1012 VSS.n1314 VSS.t1834 162.724
R1013 VSS.n1313 VSS.t1707 162.724
R1014 VSS.n1312 VSS.t1806 162.724
R1015 VSS.n1311 VSS.t1646 162.724
R1016 VSS.n1310 VSS.t457 162.724
R1017 VSS.n1261 VSS.t1859 162.724
R1018 VSS.n1260 VSS.t2122 162.724
R1019 VSS.n1259 VSS.t1671 162.724
R1020 VSS.n1258 VSS.t2462 162.724
R1021 VSS.n1257 VSS.t60 162.724
R1022 VSS.n1256 VSS.t2176 162.724
R1023 VSS.n1255 VSS.t1821 162.724
R1024 VSS.n1254 VSS.t1941 162.724
R1025 VSS.n1253 VSS.t477 162.724
R1026 VSS.n1252 VSS.t990 162.724
R1027 VSS.n1251 VSS.t116 162.724
R1028 VSS.n1250 VSS.t1525 162.724
R1029 VSS.n1249 VSS.t1274 162.724
R1030 VSS.n1248 VSS.t1640 162.724
R1031 VSS.n1247 VSS.t1036 162.724
R1032 VSS.n1246 VSS.t484 162.724
R1033 VSS.n1197 VSS.t1420 162.724
R1034 VSS.n1196 VSS.t2004 162.724
R1035 VSS.n1195 VSS.t2059 162.724
R1036 VSS.n1194 VSS.t2377 162.724
R1037 VSS.n1193 VSS.t1418 162.724
R1038 VSS.n1192 VSS.t1050 162.724
R1039 VSS.n1191 VSS.t1133 162.724
R1040 VSS.n1190 VSS.t2173 162.724
R1041 VSS.n1189 VSS.t1094 162.724
R1042 VSS.n1188 VSS.t914 162.724
R1043 VSS.n1187 VSS.t1838 162.724
R1044 VSS.n1186 VSS.t932 162.724
R1045 VSS.n1185 VSS.t488 162.724
R1046 VSS.n1184 VSS.t1350 162.724
R1047 VSS.n1183 VSS.t2283 162.724
R1048 VSS.n1182 VSS.t1063 162.724
R1049 VSS.n1133 VSS.t2343 162.724
R1050 VSS.n1132 VSS.t1919 162.724
R1051 VSS.n1131 VSS.t1766 162.724
R1052 VSS.n1130 VSS.t1256 162.724
R1053 VSS.n1129 VSS.t2261 162.724
R1054 VSS.n1128 VSS.t1558 162.724
R1055 VSS.n1127 VSS.t79 162.724
R1056 VSS.n1126 VSS.t1692 162.724
R1057 VSS.n1125 VSS.t1228 162.724
R1058 VSS.n1124 VSS.t775 162.724
R1059 VSS.n1123 VSS.t1718 162.724
R1060 VSS.n1122 VSS.t1874 162.724
R1061 VSS.n1121 VSS.t410 162.724
R1062 VSS.n1120 VSS.t1666 162.724
R1063 VSS.n1119 VSS.t868 162.724
R1064 VSS.n1118 VSS.t421 162.724
R1065 VSS.n988 VSS.t1237 162.724
R1066 VSS.n987 VSS.t382 162.724
R1067 VSS.n986 VSS.t806 162.724
R1068 VSS.n985 VSS.t1466 162.724
R1069 VSS.n984 VSS.t1276 162.724
R1070 VSS.n983 VSS.t432 162.724
R1071 VSS.n982 VSS.t1653 162.724
R1072 VSS.n981 VSS.t438 162.724
R1073 VSS.n980 VSS.t1320 162.724
R1074 VSS.n979 VSS.t2002 162.724
R1075 VSS.n978 VSS.t1259 162.724
R1076 VSS.n977 VSS.t2020 162.724
R1077 VSS.n976 VSS.t2325 162.724
R1078 VSS.n975 VSS.t861 162.724
R1079 VSS.n974 VSS.t1075 162.724
R1080 VSS.n973 VSS.t1696 162.724
R1081 VSS.n924 VSS.t1430 162.724
R1082 VSS.n923 VSS.t1752 162.724
R1083 VSS.n922 VSS.t2162 162.724
R1084 VSS.n921 VSS.t1641 162.724
R1085 VSS.n920 VSS.t89 162.724
R1086 VSS.n919 VSS.t2088 162.724
R1087 VSS.n918 VSS.t1746 162.724
R1088 VSS.n917 VSS.t1304 162.724
R1089 VSS.n916 VSS.t1791 162.724
R1090 VSS.n915 VSS.t2498 162.724
R1091 VSS.n914 VSS.t1534 162.724
R1092 VSS.n913 VSS.t235 162.724
R1093 VSS.n912 VSS.t1354 162.724
R1094 VSS.n911 VSS.t2038 162.724
R1095 VSS.n910 VSS.t953 162.724
R1096 VSS.n909 VSS.t2152 162.724
R1097 VSS.n860 VSS.t1216 162.724
R1098 VSS.n859 VSS.t1272 162.724
R1099 VSS.n858 VSS.t1841 162.724
R1100 VSS.n857 VSS.t2346 162.724
R1101 VSS.n856 VSS.t1509 162.724
R1102 VSS.n855 VSS.t1585 162.724
R1103 VSS.n854 VSS.t2148 162.724
R1104 VSS.n853 VSS.t472 162.724
R1105 VSS.n852 VSS.t2057 162.724
R1106 VSS.n851 VSS.t1185 162.724
R1107 VSS.n850 VSS.t2341 162.724
R1108 VSS.n849 VSS.t860 162.724
R1109 VSS.n848 VSS.t1794 162.724
R1110 VSS.n847 VSS.t1270 162.724
R1111 VSS.n846 VSS.t1392 162.724
R1112 VSS.n845 VSS.t2203 162.724
R1113 VSS.n796 VSS.t1290 162.724
R1114 VSS.n795 VSS.t1448 162.724
R1115 VSS.n794 VSS.t80 162.724
R1116 VSS.n793 VSS.t2195 162.724
R1117 VSS.n792 VSS.t856 162.724
R1118 VSS.n791 VSS.t1343 162.724
R1119 VSS.n790 VSS.t1830 162.724
R1120 VSS.n789 VSS.t771 162.724
R1121 VSS.n788 VSS.t1215 162.724
R1122 VSS.n787 VSS.t2262 162.724
R1123 VSS.n786 VSS.t2501 162.724
R1124 VSS.n785 VSS.t1893 162.724
R1125 VSS.n784 VSS.t2120 162.724
R1126 VSS.n783 VSS.t2110 162.724
R1127 VSS.n782 VSS.t889 162.724
R1128 VSS.n781 VSS.t2329 162.724
R1129 VSS.n700 VSS.t1403 162.724
R1130 VSS.n699 VSS.t1227 162.724
R1131 VSS.n698 VSS.t1339 162.724
R1132 VSS.n697 VSS.t1059 162.724
R1133 VSS.n696 VSS.t1096 162.724
R1134 VSS.n695 VSS.t2486 162.724
R1135 VSS.n694 VSS.t934 162.724
R1136 VSS.n693 VSS.t1912 162.724
R1137 VSS.n692 VSS.t1817 162.724
R1138 VSS.n691 VSS.t1070 162.724
R1139 VSS.n690 VSS.t854 162.724
R1140 VSS.n689 VSS.t1516 162.724
R1141 VSS.n688 VSS.t229 162.724
R1142 VSS.n687 VSS.t1845 162.724
R1143 VSS.n686 VSS.t1993 162.724
R1144 VSS.n685 VSS.t1318 162.724
R1145 VSS.n491 VSS.t2522 162.724
R1146 VSS.n490 VSS.t1402 162.724
R1147 VSS.n489 VSS.t834 162.724
R1148 VSS.n488 VSS.t1526 162.724
R1149 VSS.n487 VSS.t1358 162.724
R1150 VSS.n486 VSS.t1048 162.724
R1151 VSS.n485 VSS.t1406 162.724
R1152 VSS.n484 VSS.t2287 162.724
R1153 VSS.n483 VSS.t1851 162.724
R1154 VSS.n482 VSS.t1602 162.724
R1155 VSS.n481 VSS.t1408 162.724
R1156 VSS.n480 VSS.t881 162.724
R1157 VSS.n479 VSS.t1810 162.724
R1158 VSS.n478 VSS.t778 162.724
R1159 VSS.n477 VSS.t1179 162.724
R1160 VSS.n476 VSS.t1528 162.724
R1161 VSS.n2272 VSS.t2270 156.077
R1162 VSS.n2271 VSS.t963 156.077
R1163 VSS.n2270 VSS.t1161 156.077
R1164 VSS.n2269 VSS.t1903 156.077
R1165 VSS.n2268 VSS.t1910 156.077
R1166 VSS.n2267 VSS.t1875 156.077
R1167 VSS.n2266 VSS.t766 156.077
R1168 VSS.n2265 VSS.t2366 156.077
R1169 VSS.n2264 VSS.t2443 156.077
R1170 VSS.n2263 VSS.t2311 156.077
R1171 VSS.n2262 VSS.t2185 156.077
R1172 VSS.n2261 VSS.t2335 156.077
R1173 VSS.n2260 VSS.t896 156.077
R1174 VSS.n2259 VSS.t2452 156.077
R1175 VSS.n2258 VSS.t1965 156.077
R1176 VSS.n2257 VSS.t1191 156.077
R1177 VSS.n2176 VSS.t2309 156.077
R1178 VSS.n2175 VSS.t1459 156.077
R1179 VSS.n2174 VSS.t1139 156.077
R1180 VSS.n2173 VSS.t1719 156.077
R1181 VSS.n2172 VSS.t1617 156.077
R1182 VSS.n2171 VSS.t886 156.077
R1183 VSS.n2170 VSS.t1960 156.077
R1184 VSS.n2169 VSS.t240 156.077
R1185 VSS.n2168 VSS.t2253 156.077
R1186 VSS.n2167 VSS.t2161 156.077
R1187 VSS.n2166 VSS.t958 156.077
R1188 VSS.n2165 VSS.t1344 156.077
R1189 VSS.n2164 VSS.t1441 156.077
R1190 VSS.n2163 VSS.t878 156.077
R1191 VSS.n2162 VSS.t1870 156.077
R1192 VSS.n2161 VSS.t1078 156.077
R1193 VSS.n1950 VSS.t2011 156.077
R1194 VSS.n1949 VSS.t1296 156.077
R1195 VSS.n1948 VSS.t2496 156.077
R1196 VSS.n1947 VSS.t2351 156.077
R1197 VSS.n1946 VSS.t231 156.077
R1198 VSS.n1945 VSS.t1031 156.077
R1199 VSS.n1944 VSS.t1143 156.077
R1200 VSS.n1943 VSS.t2354 156.077
R1201 VSS.n1942 VSS.t1085 156.077
R1202 VSS.n1941 VSS.t1383 156.077
R1203 VSS.n1940 VSS.t1360 156.077
R1204 VSS.n1939 VSS.t1195 156.077
R1205 VSS.n1938 VSS.t2150 156.077
R1206 VSS.n1937 VSS.t2089 156.077
R1207 VSS.n1936 VSS.t1569 156.077
R1208 VSS.n1935 VSS.t2521 156.077
R1209 VSS.n1854 VSS.t2255 156.077
R1210 VSS.n1853 VSS.t244 156.077
R1211 VSS.n1852 VSS.t1796 156.077
R1212 VSS.n1851 VSS.t1147 156.077
R1213 VSS.n1850 VSS.t1439 156.077
R1214 VSS.n1849 VSS.t1750 156.077
R1215 VSS.n1848 VSS.t1973 156.077
R1216 VSS.n1847 VSS.t1091 156.077
R1217 VSS.n1846 VSS.t962 156.077
R1218 VSS.n1845 VSS.t2218 156.077
R1219 VSS.n1844 VSS.t1970 156.077
R1220 VSS.n1843 VSS.t115 156.077
R1221 VSS.n1842 VSS.t1363 156.077
R1222 VSS.n1841 VSS.t1450 156.077
R1223 VSS.n1840 VSS.t1715 156.077
R1224 VSS.n1839 VSS.t981 156.077
R1225 VSS.n1790 VSS.t2119 156.077
R1226 VSS.n1789 VSS.t1908 156.077
R1227 VSS.n1788 VSS.t1331 156.077
R1228 VSS.n1787 VSS.t2488 156.077
R1229 VSS.n1786 VSS.t1371 156.077
R1230 VSS.n1785 VSS.t1151 156.077
R1231 VSS.n1784 VSS.t159 156.077
R1232 VSS.n1783 VSS.t505 156.077
R1233 VSS.n1782 VSS.t1785 156.077
R1234 VSS.n1781 VSS.t1187 156.077
R1235 VSS.n1780 VSS.t1034 156.077
R1236 VSS.n1779 VSS.t497 156.077
R1237 VSS.n1778 VSS.t1258 156.077
R1238 VSS.n1777 VSS.t1894 156.077
R1239 VSS.n1776 VSS.t463 156.077
R1240 VSS.n1775 VSS.t1033 156.077
R1241 VSS.n1726 VSS.t842 156.077
R1242 VSS.n1725 VSS.t922 156.077
R1243 VSS.n1724 VSS.t2448 156.077
R1244 VSS.n1723 VSS.t467 156.077
R1245 VSS.n1722 VSS.t1802 156.077
R1246 VSS.n1721 VSS.t2485 156.077
R1247 VSS.n1720 VSS.t1163 156.077
R1248 VSS.n1719 VSS.t1545 156.077
R1249 VSS.n1718 VSS.t1315 156.077
R1250 VSS.n1717 VSS.t1453 156.077
R1251 VSS.n1716 VSS.t2052 156.077
R1252 VSS.n1715 VSS.t1975 156.077
R1253 VSS.n1714 VSS.t808 156.077
R1254 VSS.n1713 VSS.t398 156.077
R1255 VSS.n1712 VSS.t2432 156.077
R1256 VSS.n1711 VSS.t444 156.077
R1257 VSS.n1662 VSS.t1120 156.077
R1258 VSS.n1661 VSS.t894 156.077
R1259 VSS.n1660 VSS.t1346 156.077
R1260 VSS.n1659 VSS.t2181 156.077
R1261 VSS.n1658 VSS.t1100 156.077
R1262 VSS.n1657 VSS.t1041 156.077
R1263 VSS.n1656 VSS.t2278 156.077
R1264 VSS.n1655 VSS.t1622 156.077
R1265 VSS.n1654 VSS.t2503 156.077
R1266 VSS.n1653 VSS.t250 156.077
R1267 VSS.n1652 VSS.t773 156.077
R1268 VSS.n1651 VSS.t150 156.077
R1269 VSS.n1650 VSS.t1885 156.077
R1270 VSS.n1649 VSS.t1634 156.077
R1271 VSS.n1648 VSS.t2269 156.077
R1272 VSS.n1647 VSS.t2330 156.077
R1273 VSS.n1517 VSS.t809 156.077
R1274 VSS.n1516 VSS.t503 156.077
R1275 VSS.n1515 VSS.t786 156.077
R1276 VSS.n1514 VSS.t1897 156.077
R1277 VSS.n1513 VSS.t1775 156.077
R1278 VSS.n1512 VSS.t1609 156.077
R1279 VSS.n1511 VSS.t1563 156.077
R1280 VSS.n1510 VSS.t2359 156.077
R1281 VSS.n1509 VSS.t66 156.077
R1282 VSS.n1508 VSS.t1722 156.077
R1283 VSS.n1507 VSS.t999 156.077
R1284 VSS.n1506 VSS.t1765 156.077
R1285 VSS.n1505 VSS.t447 156.077
R1286 VSS.n1504 VSS.t1531 156.077
R1287 VSS.n1503 VSS.t1477 156.077
R1288 VSS.n1502 VSS.t253 156.077
R1289 VSS.n1453 VSS.t2163 156.077
R1290 VSS.n1452 VSS.t1113 156.077
R1291 VSS.n1451 VSS.t1782 156.077
R1292 VSS.n1450 VSS.t507 156.077
R1293 VSS.n1449 VSS.t816 156.077
R1294 VSS.n1448 VSS.t1582 156.077
R1295 VSS.n1447 VSS.t1167 156.077
R1296 VSS.n1446 VSS.t2211 156.077
R1297 VSS.n1445 VSS.t942 156.077
R1298 VSS.n1444 VSS.t2136 156.077
R1299 VSS.n1443 VSS.t2045 156.077
R1300 VSS.n1442 VSS.t1962 156.077
R1301 VSS.n1441 VSS.t955 156.077
R1302 VSS.n1440 VSS.t1201 156.077
R1303 VSS.n1439 VSS.t2079 156.077
R1304 VSS.n1438 VSS.t916 156.077
R1305 VSS.n1389 VSS.t417 156.077
R1306 VSS.n1388 VSS.t1038 156.077
R1307 VSS.n1387 VSS.t2092 156.077
R1308 VSS.n1386 VSS.t1819 156.077
R1309 VSS.n1385 VSS.t1000 156.077
R1310 VSS.n1384 VSS.t2124 156.077
R1311 VSS.n1383 VSS.t1482 156.077
R1312 VSS.n1382 VSS.t249 156.077
R1313 VSS.n1381 VSS.t2342 156.077
R1314 VSS.n1380 VSS.t2147 156.077
R1315 VSS.n1379 VSS.t1789 156.077
R1316 VSS.n1378 VSS.t2105 156.077
R1317 VSS.n1377 VSS.t2468 156.077
R1318 VSS.n1376 VSS.t1442 156.077
R1319 VSS.n1375 VSS.t1590 156.077
R1320 VSS.n1374 VSS.t1056 156.077
R1321 VSS.n1325 VSS.t925 156.077
R1322 VSS.n1324 VSS.t2238 156.077
R1323 VSS.n1323 VSS.t1881 156.077
R1324 VSS.n1322 VSS.t1455 156.077
R1325 VSS.n1321 VSS.t1382 156.077
R1326 VSS.n1320 VSS.t976 156.077
R1327 VSS.n1319 VSS.t1175 156.077
R1328 VSS.n1318 VSS.t50 156.077
R1329 VSS.n1317 VSS.t1188 156.077
R1330 VSS.n1316 VSS.t1551 156.077
R1331 VSS.n1315 VSS.t439 156.077
R1332 VSS.n1314 VSS.t1835 156.077
R1333 VSS.n1313 VSS.t1708 156.077
R1334 VSS.n1312 VSS.t1805 156.077
R1335 VSS.n1311 VSS.t433 156.077
R1336 VSS.n1310 VSS.t456 156.077
R1337 VSS.n1261 VSS.t1860 156.077
R1338 VSS.n1260 VSS.t1060 156.077
R1339 VSS.n1259 VSS.t1670 156.077
R1340 VSS.n1258 VSS.t2472 156.077
R1341 VSS.n1257 VSS.t65 156.077
R1342 VSS.n1256 VSS.t2339 156.077
R1343 VSS.n1255 VSS.t1347 156.077
R1344 VSS.n1254 VSS.t1940 156.077
R1345 VSS.n1253 VSS.t476 156.077
R1346 VSS.n1252 VSS.t989 156.077
R1347 VSS.n1251 VSS.t109 156.077
R1348 VSS.n1250 VSS.t1524 156.077
R1349 VSS.n1249 VSS.t1273 156.077
R1350 VSS.n1248 VSS.t1639 156.077
R1351 VSS.n1247 VSS.t1037 156.077
R1352 VSS.n1246 VSS.t483 156.077
R1353 VSS.n1197 VSS.t1421 156.077
R1354 VSS.n1196 VSS.t1278 156.077
R1355 VSS.n1195 VSS.t2128 156.077
R1356 VSS.n1194 VSS.t2378 156.077
R1357 VSS.n1193 VSS.t1419 156.077
R1358 VSS.n1192 VSS.t1049 156.077
R1359 VSS.n1191 VSS.t1132 156.077
R1360 VSS.n1190 VSS.t2367 156.077
R1361 VSS.n1189 VSS.t1095 156.077
R1362 VSS.n1188 VSS.t913 156.077
R1363 VSS.n1187 VSS.t1848 156.077
R1364 VSS.n1186 VSS.t931 156.077
R1365 VSS.n1185 VSS.t1781 156.077
R1366 VSS.n1184 VSS.t1349 156.077
R1367 VSS.n1183 VSS.t2284 156.077
R1368 VSS.n1182 VSS.t1062 156.077
R1369 VSS.n1133 VSS.t2338 156.077
R1370 VSS.n1132 VSS.t1918 156.077
R1371 VSS.n1131 VSS.t1767 156.077
R1372 VSS.n1130 VSS.t1255 156.077
R1373 VSS.n1129 VSS.t2201 156.077
R1374 VSS.n1128 VSS.t1557 156.077
R1375 VSS.n1127 VSS.t78 156.077
R1376 VSS.n1126 VSS.t838 156.077
R1377 VSS.n1125 VSS.t1229 156.077
R1378 VSS.n1124 VSS.t774 156.077
R1379 VSS.n1123 VSS.t1717 156.077
R1380 VSS.n1122 VSS.t1832 156.077
R1381 VSS.n1121 VSS.t411 156.077
R1382 VSS.n1120 VSS.t1665 156.077
R1383 VSS.n1119 VSS.t867 156.077
R1384 VSS.n1118 VSS.t420 156.077
R1385 VSS.n988 VSS.t1238 156.077
R1386 VSS.n987 VSS.t404 156.077
R1387 VSS.n986 VSS.t805 156.077
R1388 VSS.n985 VSS.t1465 156.077
R1389 VSS.n984 VSS.t1277 156.077
R1390 VSS.n983 VSS.t431 156.077
R1391 VSS.n982 VSS.t2280 156.077
R1392 VSS.n981 VSS.t440 156.077
R1393 VSS.n980 VSS.t1321 156.077
R1394 VSS.n979 VSS.t2003 156.077
R1395 VSS.n978 VSS.t1275 156.077
R1396 VSS.n977 VSS.t2019 156.077
R1397 VSS.n976 VSS.t2266 156.077
R1398 VSS.n975 VSS.t1566 156.077
R1399 VSS.n974 VSS.t940 156.077
R1400 VSS.n973 VSS.t1695 156.077
R1401 VSS.n924 VSS.t1431 156.077
R1402 VSS.n923 VSS.t1417 156.077
R1403 VSS.n922 VSS.t2235 156.077
R1404 VSS.n921 VSS.t1647 156.077
R1405 VSS.n920 VSS.t83 156.077
R1406 VSS.n919 VSS.t2087 156.077
R1407 VSS.n918 VSS.t1747 156.077
R1408 VSS.n917 VSS.t1303 156.077
R1409 VSS.n916 VSS.t1790 156.077
R1410 VSS.n915 VSS.t2497 156.077
R1411 VSS.n914 VSS.t1535 156.077
R1412 VSS.n913 VSS.t241 156.077
R1413 VSS.n912 VSS.t1355 156.077
R1414 VSS.n911 VSS.t2037 156.077
R1415 VSS.n910 VSS.t952 156.077
R1416 VSS.n909 VSS.t2276 156.077
R1417 VSS.n860 VSS.t1217 156.077
R1418 VSS.n859 VSS.t1271 156.077
R1419 VSS.n858 VSS.t1840 156.077
R1420 VSS.n857 VSS.t2345 156.077
R1421 VSS.n856 VSS.t1180 156.077
R1422 VSS.n855 VSS.t1584 156.077
R1423 VSS.n854 VSS.t1325 156.077
R1424 VSS.n853 VSS.t473 156.077
R1425 VSS.n852 VSS.t2058 156.077
R1426 VSS.n851 VSS.t1184 156.077
R1427 VSS.n850 VSS.t2340 156.077
R1428 VSS.n849 VSS.t2332 156.077
R1429 VSS.n848 VSS.t1795 156.077
R1430 VSS.n847 VSS.t1269 156.077
R1431 VSS.n846 VSS.t1391 156.077
R1432 VSS.n845 VSS.t2202 156.077
R1433 VSS.n796 VSS.t1291 156.077
R1434 VSS.n795 VSS.t1447 156.077
R1435 VSS.n794 VSS.t81 156.077
R1436 VSS.n793 VSS.t2196 156.077
R1437 VSS.n792 VSS.t857 156.077
R1438 VSS.n791 VSS.t1342 156.077
R1439 VSS.n790 VSS.t1833 156.077
R1440 VSS.n789 VSS.t770 156.077
R1441 VSS.n788 VSS.t1214 156.077
R1442 VSS.n787 VSS.t2440 156.077
R1443 VSS.n786 VSS.t2500 156.077
R1444 VSS.n785 VSS.t1892 156.077
R1445 VSS.n784 VSS.t2121 156.077
R1446 VSS.n783 VSS.t2109 156.077
R1447 VSS.n782 VSS.t888 156.077
R1448 VSS.n781 VSS.t2260 156.077
R1449 VSS.n700 VSS.t1404 156.077
R1450 VSS.n699 VSS.t1226 156.077
R1451 VSS.n698 VSS.t1338 156.077
R1452 VSS.n697 VSS.t1648 156.077
R1453 VSS.n696 VSS.t1097 156.077
R1454 VSS.n695 VSS.t2480 156.077
R1455 VSS.n694 VSS.t933 156.077
R1456 VSS.n693 VSS.t1911 156.077
R1457 VSS.n692 VSS.t1818 156.077
R1458 VSS.n691 VSS.t1072 156.077
R1459 VSS.n690 VSS.t480 156.077
R1460 VSS.n689 VSS.t1515 156.077
R1461 VSS.n688 VSS.t114 156.077
R1462 VSS.n687 VSS.t1844 156.077
R1463 VSS.n686 VSS.t1992 156.077
R1464 VSS.n685 VSS.t1319 156.077
R1465 VSS.n573 VSS.t2171 156.077
R1466 VSS.n576 VSS.t64 156.077
R1467 VSS.n618 VSS.t2013 156.077
R1468 VSS.n1610 VSS.t487 156.077
R1469 VSS.n2093 VSS.t1689 156.077
R1470 VSS.n1081 VSS.t1549 156.077
R1471 VSS.n615 VSS.t1571 156.077
R1472 VSS.n1607 VSS.t2183 156.077
R1473 VSS.n2089 VSS.t2154 156.077
R1474 VSS.n1078 VSS.t2094 156.077
R1475 VSS.n612 VSS.t1374 156.077
R1476 VSS.n1604 VSS.t2520 156.077
R1477 VSS.n2085 VSS.t1742 156.077
R1478 VSS.n1075 VSS.t1854 156.077
R1479 VSS.n609 VSS.t1861 156.077
R1480 VSS.n1601 VSS.t2036 156.077
R1481 VSS.n2081 VSS.t2248 156.077
R1482 VSS.n1072 VSS.t1137 156.077
R1483 VSS.n606 VSS.t1105 156.077
R1484 VSS.n1598 VSS.t94 156.077
R1485 VSS.n2077 VSS.t2510 156.077
R1486 VSS.n1069 VSS.t462 156.077
R1487 VSS.n603 VSS.t1323 156.077
R1488 VSS.n1595 VSS.t2527 156.077
R1489 VSS.n2073 VSS.t1457 156.077
R1490 VSS.n1066 VSS.t817 156.077
R1491 VSS.n600 VSS.t898 156.077
R1492 VSS.n1592 VSS.t1434 156.077
R1493 VSS.n2069 VSS.t2138 156.077
R1494 VSS.n1063 VSS.t2293 156.077
R1495 VSS.n597 VSS.t2328 156.077
R1496 VSS.n1589 VSS.t1703 156.077
R1497 VSS.n2065 VSS.t924 156.077
R1498 VSS.n1060 VSS.t929 156.077
R1499 VSS.n594 VSS.t2484 156.077
R1500 VSS.n1586 VSS.t2108 156.077
R1501 VSS.n2061 VSS.t1604 156.077
R1502 VSS.n1057 VSS.t980 156.077
R1503 VSS.n591 VSS.t1054 156.077
R1504 VSS.n1583 VSS.t30 156.077
R1505 VSS.n2057 VSS.t57 156.077
R1506 VSS.n1054 VSS.t1480 156.077
R1507 VSS.n588 VSS.t2070 156.077
R1508 VSS.n1580 VSS.t1288 156.077
R1509 VSS.n2053 VSS.t392 156.077
R1510 VSS.n1051 VSS.t871 156.077
R1511 VSS.n585 VSS.t1111 156.077
R1512 VSS.n1577 VSS.t1738 156.077
R1513 VSS.n2049 VSS.t2190 156.077
R1514 VSS.n1048 VSS.t2251 156.077
R1515 VSS.n582 VSS.t1093 156.077
R1516 VSS.n1574 VSS.t879 156.077
R1517 VSS.n2045 VSS.t1995 156.077
R1518 VSS.n1045 VSS.t2028 156.077
R1519 VSS.n579 VSS.t1127 156.077
R1520 VSS.n1571 VSS.t997 156.077
R1521 VSS.n2041 VSS.t46 156.077
R1522 VSS.n1042 VSS.t1886 156.077
R1523 VSS.n1038 VSS.t768 156.077
R1524 VSS.n1113 VSS.t1284 156.077
R1525 VSS.n2037 VSS.t1677 156.077
R1526 VSS.n1568 VSS.t850 156.077
R1527 VSS.n1644 VSS.t1899 156.077
R1528 VSS.n2033 VSS.t2265 156.077
R1529 VSS.n491 VSS.t2502 156.077
R1530 VSS.n490 VSS.t1401 156.077
R1531 VSS.n489 VSS.t833 156.077
R1532 VSS.n488 VSS.t1487 156.077
R1533 VSS.n487 VSS.t1359 156.077
R1534 VSS.n486 VSS.t1047 156.077
R1535 VSS.n485 VSS.t1405 156.077
R1536 VSS.n484 VSS.t2286 156.077
R1537 VSS.n483 VSS.t1852 156.077
R1538 VSS.n482 VSS.t1601 156.077
R1539 VSS.n481 VSS.t1407 156.077
R1540 VSS.n480 VSS.t1967 156.077
R1541 VSS.n479 VSS.t1811 156.077
R1542 VSS.n478 VSS.t777 156.077
R1543 VSS.n477 VSS.t1178 156.077
R1544 VSS.n476 VSS.t1527 156.077
R1545 VSS.n2221 VSS.t1194 154.891
R1546 VSS.n2218 VSS.t1964 154.891
R1547 VSS.n2215 VSS.t2427 154.891
R1548 VSS.n2212 VSS.t1379 154.891
R1549 VSS.n2209 VSS.t2174 154.891
R1550 VSS.n2206 VSS.t2180 154.891
R1551 VSS.n2203 VSS.t2424 154.891
R1552 VSS.n2200 VSS.t2430 154.891
R1553 VSS.n2197 VSS.t2371 154.891
R1554 VSS.n2194 VSS.t1997 154.891
R1555 VSS.n2191 VSS.t1864 154.891
R1556 VSS.n2188 VSS.t1197 154.891
R1557 VSS.n2185 VSS.t1706 154.891
R1558 VSS.n2182 VSS.t2450 154.891
R1559 VSS.n2179 VSS.t1917 154.891
R1560 VSS.n2177 VSS.t2364 154.891
R1561 VSS.n1995 VSS.t2322 154.891
R1562 VSS.n1992 VSS.t1337 154.891
R1563 VSS.n1989 VSS.t1773 154.891
R1564 VSS.n1986 VSS.t1605 154.891
R1565 VSS.n1983 VSS.t2347 154.891
R1566 VSS.n1980 VSS.t391 154.891
R1567 VSS.n1977 VSS.t2363 154.891
R1568 VSS.n1974 VSS.t1043 154.891
R1569 VSS.n1971 VSS.t1110 154.891
R1570 VSS.n1968 VSS.t1148 154.891
R1571 VSS.n1965 VSS.t1888 154.891
R1572 VSS.n1962 VSS.t2511 154.891
R1573 VSS.n1959 VSS.t2250 154.891
R1574 VSS.n1956 VSS.t1932 154.891
R1575 VSS.n1953 VSS.t969 154.891
R1576 VSS.n1951 VSS.t1741 154.891
R1577 VSS.n1899 VSS.t2490 154.891
R1578 VSS.n1896 VSS.t1568 154.891
R1579 VSS.n1893 VSS.t1779 154.891
R1580 VSS.n1890 VSS.t2146 154.891
R1581 VSS.n1887 VSS.t1182 154.891
R1582 VSS.n1884 VSS.t2294 154.891
R1583 VSS.n1881 VSS.t1685 154.891
R1584 VSS.n1878 VSS.t1134 154.891
R1585 VSS.n1875 VSS.t1824 154.891
R1586 VSS.n1872 VSS.t1592 154.891
R1587 VSS.n1869 VSS.t1028 154.891
R1588 VSS.n1866 VSS.t104 154.891
R1589 VSS.n1863 VSS.t2350 154.891
R1590 VSS.n1860 VSS.t2246 154.891
R1591 VSS.n1857 VSS.t2010 154.891
R1592 VSS.n1855 VSS.t1611 154.891
R1593 VSS.n1835 VSS.t2047 154.891
R1594 VSS.n1832 VSS.t1608 154.891
R1595 VSS.n1829 VSS.t1116 154.891
R1596 VSS.n1826 VSS.t1365 154.891
R1597 VSS.n1823 VSS.t232 154.891
R1598 VSS.n1820 VSS.t2055 154.891
R1599 VSS.n1817 VSS.t2213 154.891
R1600 VSS.n1814 VSS.t1506 154.891
R1601 VSS.n1811 VSS.t1199 154.891
R1602 VSS.n1808 VSS.t1771 154.891
R1603 VSS.n1805 VSS.t1710 154.891
R1604 VSS.n1802 VSS.t1436 154.891
R1605 VSS.n1799 VSS.t1006 154.891
R1606 VSS.n1796 VSS.t1645 154.891
R1607 VSS.n1793 VSS.t245 154.891
R1608 VSS.n1791 VSS.t2257 154.891
R1609 VSS.n1771 VSS.t1702 154.891
R1610 VSS.n1768 VSS.t2240 154.891
R1611 VSS.n1765 VSS.t1287 154.891
R1612 VSS.n1762 VSS.t2023 154.891
R1613 VSS.n1759 VSS.t1546 154.891
R1614 VSS.n1756 VSS.t1598 154.891
R1615 VSS.n1753 VSS.t1508 154.891
R1616 VSS.n1750 VSS.t482 154.891
R1617 VSS.n1747 VSS.t1620 154.891
R1618 VSS.n1744 VSS.t67 154.891
R1619 VSS.n1741 VSS.t1261 154.891
R1620 VSS.n1738 VSS.t1739 154.891
R1621 VSS.n1735 VSS.t153 154.891
R1622 VSS.n1732 VSS.t1334 154.891
R1623 VSS.n1729 VSS.t1263 154.891
R1624 VSS.n1727 VSS.t491 154.891
R1625 VSS.n1707 VSS.t1057 154.891
R1626 VSS.n1704 VSS.t85 154.891
R1627 VSS.n1701 VSS.t1533 154.891
R1628 VSS.n1698 VSS.t1472 154.891
R1629 VSS.n1695 VSS.t848 154.891
R1630 VSS.n1692 VSS.t2051 154.891
R1631 VSS.n1689 VSS.t1451 154.891
R1632 VSS.n1686 VSS.t1166 154.891
R1633 VSS.n1683 VSS.t1544 154.891
R1634 VSS.n1680 VSS.t2083 154.891
R1635 VSS.n1677 VSS.t2327 154.891
R1636 VSS.n1674 VSS.t2323 154.891
R1637 VSS.n1671 VSS.t464 154.891
R1638 VSS.n1668 VSS.t902 154.891
R1639 VSS.n1665 VSS.t1829 154.891
R1640 VSS.n1663 VSS.t436 154.891
R1641 VSS.n1562 VSS.t1589 154.891
R1642 VSS.n1559 VSS.t1539 154.891
R1643 VSS.n1556 VSS.t994 154.891
R1644 VSS.n1553 VSS.t1177 154.891
R1645 VSS.n1550 VSS.t1882 154.891
R1646 VSS.n1547 VSS.t1628 154.891
R1647 VSS.n1544 VSS.t44 154.891
R1648 VSS.n1541 VSS.t2299 154.891
R1649 VSS.n1538 VSS.t2001 154.891
R1650 VSS.n1535 VSS.t791 154.891
R1651 VSS.n1532 VSS.t2473 154.891
R1652 VSS.n1529 VSS.t2104 154.891
R1653 VSS.n1526 VSS.t1873 154.891
R1654 VSS.n1523 VSS.t2518 154.891
R1655 VSS.n1520 VSS.t2188 154.891
R1656 VSS.n1518 VSS.t1686 154.891
R1657 VSS.n1498 VSS.t394 154.891
R1658 VSS.n1495 VSS.t1836 154.891
R1659 VSS.n1492 VSS.t1553 154.891
R1660 VSS.n1489 VSS.t452 154.891
R1661 VSS.n1486 VSS.t1725 154.891
R1662 VSS.n1483 VSS.t1986 154.891
R1663 VSS.n1480 VSS.t1820 154.891
R1664 VSS.n1477 VSS.t2417 154.891
R1665 VSS.n1474 VSS.t55 154.891
R1666 VSS.n1471 VSS.t1561 154.891
R1667 VSS.n1468 VSS.t1799 154.891
R1668 VSS.n1465 VSS.t1029 154.891
R1669 VSS.n1462 VSS.t1456 154.891
R1670 VSS.n1459 VSS.t793 154.891
R1671 VSS.n1456 VSS.t2331 154.891
R1672 VSS.n1454 VSS.t2061 154.891
R1673 VSS.n1434 VSS.t1697 154.891
R1674 VSS.n1431 VSS.t1190 154.891
R1675 VSS.n1428 VSS.t1203 154.891
R1676 VSS.n1425 VSS.t1680 154.891
R1677 VSS.n1422 VSS.t1298 154.891
R1678 VSS.n1419 VSS.t2074 154.891
R1679 VSS.n1416 VSS.t876 154.891
R1680 VSS.n1413 VSS.t1842 154.891
R1681 VSS.n1410 VSS.t2217 154.891
R1682 VSS.n1407 VSS.t1687 154.891
R1683 VSS.n1404 VSS.t966 154.891
R1684 VSS.n1401 VSS.t1869 154.891
R1685 VSS.n1398 VSS.t1613 154.891
R1686 VSS.n1395 VSS.t2256 154.891
R1687 VSS.n1392 VSS.t1429 154.891
R1688 VSS.n1390 VSS.t2307 154.891
R1689 VSS.n1370 VSS.t1847 154.891
R1690 VSS.n1367 VSS.t1594 154.891
R1691 VSS.n1364 VSS.t1826 154.891
R1692 VSS.n1361 VSS.t2478 154.891
R1693 VSS.n1358 VSS.t1015 154.891
R1694 VSS.n1355 VSS.t1649 154.891
R1695 VSS.n1352 VSS.t1311 154.891
R1696 VSS.n1349 VSS.t407 154.891
R1697 VSS.n1346 VSS.t228 154.891
R1698 VSS.n1343 VSS.t499 154.891
R1699 VSS.n1340 VSS.t434 154.891
R1700 VSS.n1337 VSS.t1076 154.891
R1701 VSS.n1334 VSS.t424 154.891
R1702 VSS.n1331 VSS.t1142 154.891
R1703 VSS.n1328 VSS.t2170 154.891
R1704 VSS.n1326 VSS.t2142 154.891
R1705 VSS.n1306 VSS.t468 154.891
R1706 VSS.n1303 VSS.t974 154.891
R1707 VSS.n1300 VSS.t837 154.891
R1708 VSS.n1297 VSS.t2040 154.891
R1709 VSS.n1294 VSS.t1425 154.891
R1710 VSS.n1291 VSS.t1317 154.891
R1711 VSS.n1288 VSS.t1651 154.891
R1712 VSS.n1285 VSS.t1510 154.891
R1713 VSS.n1282 VSS.t1793 154.891
R1714 VSS.n1279 VSS.t1683 154.891
R1715 VSS.n1276 VSS.t2065 154.891
R1716 VSS.n1273 VSS.t1808 154.891
R1717 VSS.n1270 VSS.t2050 154.891
R1718 VSS.n1267 VSS.t1219 154.891
R1719 VSS.n1264 VSS.t1968 154.891
R1720 VSS.n1262 VSS.t1637 154.891
R1721 VSS.n1242 VSS.t471 154.891
R1722 VSS.n1239 VSS.t2144 154.891
R1723 VSS.n1236 VSS.t2156 154.891
R1724 VSS.n1233 VSS.t1769 154.891
R1725 VSS.n1230 VSS.t2081 154.891
R1726 VSS.n1227 VSS.t388 154.891
R1727 VSS.n1224 VSS.t426 154.891
R1728 VSS.n1221 VSS.t855 154.891
R1729 VSS.n1218 VSS.t1943 154.891
R1730 VSS.n1215 VSS.t1330 154.891
R1731 VSS.n1212 VSS.t1959 154.891
R1732 VSS.n1209 VSS.t47 154.891
R1733 VSS.n1206 VSS.t2475 154.891
R1734 VSS.n1203 VSS.t1667 154.891
R1735 VSS.n1200 VSS.t1101 154.891
R1736 VSS.n1198 VSS.t2076 154.891
R1737 VSS.n1178 VSS.t1675 154.891
R1738 VSS.n1175 VSS.t2279 154.891
R1739 VSS.n1172 VSS.t1556 154.891
R1740 VSS.n1169 VSS.t1326 154.891
R1741 VSS.n1166 VSS.t904 154.891
R1742 VSS.n1163 VSS.t1839 154.891
R1743 VSS.n1160 VSS.t872 154.891
R1744 VSS.n1157 VSS.t1071 154.891
R1745 VSS.n1154 VSS.t1517 154.891
R1746 VSS.n1151 VSS.t1335 154.891
R1747 VSS.n1148 VSS.t1476 154.891
R1748 VSS.n1145 VSS.t502 154.891
R1749 VSS.n1142 VSS.t2375 154.891
R1750 VSS.n1139 VSS.t891 154.891
R1751 VSS.n1136 VSS.t823 154.891
R1752 VSS.n1134 VSS.t852 154.891
R1753 VSS.n1033 VSS.t1136 154.891
R1754 VSS.n1030 VSS.t1373 154.891
R1755 VSS.n1027 VSS.t798 154.891
R1756 VSS.n1024 VSS.t1233 154.891
R1757 VSS.n1021 VSS.t2244 154.891
R1758 VSS.n1018 VSS.t1003 154.891
R1759 VSS.n1015 VSS.t2008 154.891
R1760 VSS.n1012 VSS.t1357 154.891
R1761 VSS.n1009 VSS.t928 154.891
R1762 VSS.n1006 VSS.t926 154.891
R1763 VSS.n1003 VSS.t1921 154.891
R1764 VSS.n1000 VSS.t804 154.891
R1765 VSS.n997 VSS.t1736 154.891
R1766 VSS.n994 VSS.t1253 154.891
R1767 VSS.n991 VSS.t2127 154.891
R1768 VSS.n989 VSS.t1411 154.891
R1769 VSS.n969 VSS.t947 154.891
R1770 VSS.n966 VSS.t2077 154.891
R1771 VSS.n963 VSS.t1756 154.891
R1772 VSS.n960 VSS.t2508 154.891
R1773 VSS.n957 VSS.t2021 154.891
R1774 VSS.n954 VSS.t1822 154.891
R1775 VSS.n951 VSS.t2005 154.891
R1776 VSS.n948 VSS.t1906 154.891
R1777 VSS.n945 VSS.t1514 154.891
R1778 VSS.n942 VSS.t475 154.891
R1779 VSS.n939 VSS.t1489 154.891
R1780 VSS.n936 VSS.t1559 154.891
R1781 VSS.n933 VSS.t1987 154.891
R1782 VSS.n930 VSS.t409 154.891
R1783 VSS.n927 VSS.t242 154.891
R1784 VSS.n925 VSS.t1206 154.891
R1785 VSS.n905 VSS.t2273 154.891
R1786 VSS.n902 VSS.t1804 154.891
R1787 VSS.n899 VSS.t1914 154.891
R1788 VSS.n896 VSS.t821 154.891
R1789 VSS.n893 VSS.t1555 154.891
R1790 VSS.n890 VSS.t2449 154.891
R1791 VSS.n887 VSS.t2495 154.891
R1792 VSS.n884 VSS.t2053 154.891
R1793 VSS.n881 VSS.t1306 154.891
R1794 VSS.n878 VSS.t1051 154.891
R1795 VSS.n875 VSS.t1146 154.891
R1796 VSS.n872 VSS.t90 154.891
R1797 VSS.n869 VSS.t479 154.891
R1798 VSS.n866 VSS.t2310 154.891
R1799 VSS.n863 VSS.t1005 154.891
R1800 VSS.n861 VSS.t1089 154.891
R1801 VSS.n841 VSS.t2206 154.891
R1802 VSS.n838 VSS.t1393 154.891
R1803 VSS.n835 VSS.t1446 154.891
R1804 VSS.n832 VSS.t1991 154.891
R1805 VSS.n829 VSS.t2243 154.891
R1806 VSS.n826 VSS.t261 154.891
R1807 VSS.n823 VSS.t2421 154.891
R1808 VSS.n820 VSS.t1587 154.891
R1809 VSS.n817 VSS.t450 154.891
R1810 VSS.n814 VSS.t1657 154.891
R1811 VSS.n811 VSS.t2114 154.891
R1812 VSS.n808 VSS.t1933 154.891
R1813 VSS.n805 VSS.t2334 154.891
R1814 VSS.n802 VSS.t1850 154.891
R1815 VSS.n799 VSS.t1200 154.891
R1816 VSS.n797 VSS.t1626 154.891
R1817 VSS.n745 VSS.t2471 154.891
R1818 VSS.n742 VSS.t870 154.891
R1819 VSS.n739 VSS.t1990 154.891
R1820 VSS.n736 VSS.t1242 154.891
R1821 VSS.n733 VSS.t1890 154.891
R1822 VSS.n730 VSS.t2369 154.891
R1823 VSS.n727 VSS.t2447 154.891
R1824 VSS.n724 VSS.t1470 154.891
R1825 VSS.n721 VSS.t1749 154.891
R1826 VSS.n718 VSS.t1630 154.891
R1827 VSS.n715 VSS.t789 154.891
R1828 VSS.n712 VSS.t2297 154.891
R1829 VSS.n709 VSS.t2461 154.891
R1830 VSS.n706 VSS.t2358 154.891
R1831 VSS.n703 VSS.t413 154.891
R1832 VSS.n701 VSS.t1868 154.891
R1833 VSS.n574 VSS.t1730 154.891
R1834 VSS.n577 VSS.t1468 154.891
R1835 VSS.n580 VSS.t1414 154.891
R1836 VSS.n583 VSS.t386 154.891
R1837 VSS.n586 VSS.t1073 154.891
R1838 VSS.n589 VSS.t858 154.891
R1839 VSS.n592 VSS.t1090 154.891
R1840 VSS.n595 VSS.t1328 154.891
R1841 VSS.n598 VSS.t1957 154.891
R1842 VSS.n601 VSS.t935 154.891
R1843 VSS.n604 VSS.t2463 154.891
R1844 VSS.n607 VSS.t2157 154.891
R1845 VSS.n610 VSS.t1102 154.891
R1846 VSS.n613 VSS.t1266 154.891
R1847 VSS.n616 VSS.t1896 154.891
R1848 VSS.n619 VSS.t2026 154.891
R1849 VSS.n2094 VSS.t2205 154.891
R1850 VSS.n1039 VSS.t1433 154.891
R1851 VSS.n1040 VSS.t1754 154.891
R1852 VSS.n1043 VSS.t1662 154.891
R1853 VSS.n1046 VSS.t1513 154.891
R1854 VSS.n1049 VSS.t813 154.891
R1855 VSS.n1052 VSS.t1377 154.891
R1856 VSS.n1055 VSS.t1068 154.891
R1857 VSS.n1058 VSS.t2032 154.891
R1858 VSS.n1061 VSS.t2063 154.891
R1859 VSS.n1064 VSS.t1125 154.891
R1860 VSS.n1067 VSS.t1745 154.891
R1861 VSS.n1070 VSS.t2303 154.891
R1862 VSS.n1073 VSS.t419 154.891
R1863 VSS.n1076 VSS.t1797 154.891
R1864 VSS.n1079 VSS.t2112 154.891
R1865 VSS.n1082 VSS.t1976 154.891
R1866 VSS.n1566 VSS.t2482 154.891
R1867 VSS.n1569 VSS.t1250 154.891
R1868 VSS.n1572 VSS.t1295 154.891
R1869 VSS.n1575 VSS.t944 154.891
R1870 VSS.n1578 VSS.t1131 154.891
R1871 VSS.n1581 VSS.t1220 154.891
R1872 VSS.n1584 VSS.t252 154.891
R1873 VSS.n1587 VSS.t2282 154.891
R1874 VSS.n1590 VSS.t1623 154.891
R1875 VSS.n1593 VSS.t2487 154.891
R1876 VSS.n1596 VSS.t1014 154.891
R1877 VSS.n1599 VSS.t1086 154.891
R1878 VSS.n1602 VSS.t1734 154.891
R1879 VSS.n1605 VSS.t1348 154.891
R1880 VSS.n1608 VSS.t492 154.891
R1881 VSS.n1611 VSS.t1119 154.891
R1882 VSS.n2034 VSS.t912 154.891
R1883 VSS.n2038 VSS.t1758 154.891
R1884 VSS.n2042 VSS.t1463 154.891
R1885 VSS.n2046 VSS.t459 154.891
R1886 VSS.n2050 VSS.t1654 154.891
R1887 VSS.n2054 VSS.t960 154.891
R1888 VSS.n2058 VSS.t2182 154.891
R1889 VSS.n2062 VSS.t236 154.891
R1890 VSS.n2066 VSS.t108 154.891
R1891 VSS.n2070 VSS.t1632 154.891
R1892 VSS.n2074 VSS.t776 154.891
R1893 VSS.n2078 VSS.t1618 154.891
R1894 VSS.n2082 VSS.t1723 154.891
R1895 VSS.n2086 VSS.t2086 154.891
R1896 VSS.n2090 VSS.t2214 154.891
R1897 VSS.n536 VSS.t2167 154.891
R1898 VSS.n533 VSS.t61 154.891
R1899 VSS.n530 VSS.t1523 154.891
R1900 VSS.n527 VSS.t1519 154.891
R1901 VSS.n524 VSS.t945 154.891
R1902 VSS.n521 VSS.t1727 154.891
R1903 VSS.n518 VSS.t1052 154.891
R1904 VSS.n515 VSS.t2429 154.891
R1905 VSS.n512 VSS.t2441 154.891
R1906 VSS.n509 VSS.t1595 154.891
R1907 VSS.n506 VSS.t1322 154.891
R1908 VSS.n503 VSS.t1711 154.891
R1909 VSS.n500 VSS.t441 154.891
R1910 VSS.n497 VSS.t1308 154.891
R1911 VSS.n494 VSS.t796 154.891
R1912 VSS.n492 VSS.t1231 154.891
R1913 VSS.n442 VSS.t1292 154.891
R1914 VSS.n440 VSS.t1117 154.891
R1915 VSS.n438 VSS.t1635 154.891
R1916 VSS.n436 VSS.t840 154.891
R1917 VSS.n434 VSS.t1776 154.891
R1918 VSS.n432 VSS.t795 154.891
R1919 VSS.n430 VSS.t1389 154.891
R1920 VSS.n428 VSS.t1351 154.891
R1921 VSS.n426 VSS.t2492 154.891
R1922 VSS.n424 VSS.t415 154.891
R1923 VSS.n422 VSS.t1279 154.891
R1924 VSS.n420 VSS.t1239 154.891
R1925 VSS.n418 VSS.t920 154.891
R1926 VSS.n416 VSS.t1672 154.891
R1927 VSS.n414 VSS.t1170 154.891
R1928 VSS.n413 VSS.t2285 154.891
R1929 VSS.n2129 VSS.t719 154.248
R1930 VSS.n653 VSS.t725 154.248
R1931 VSS.n2225 VSS.t596 154.243
R1932 VSS.n1999 VSS.t738 154.243
R1933 VSS.n1903 VSS.t550 154.243
R1934 VSS.n749 VSS.t552 154.243
R1935 VSS.n540 VSS.t711 154.243
R1936 VSS.n444 VSS.t586 154.243
R1937 VSS.n2241 VSS.t542 154.228
R1938 VSS.n2145 VSS.t702 154.228
R1939 VSS.n2015 VSS.t724 154.228
R1940 VSS.n1919 VSS.t541 154.228
R1941 VSS.n765 VSS.t645 154.228
R1942 VSS.n669 VSS.t560 154.228
R1943 VSS.n556 VSS.t546 154.228
R1944 VSS.n460 VSS.t674 154.228
R1945 VSS.n2255 VSS.t563 149.249
R1946 VSS.n2254 VSS.t689 149.249
R1947 VSS.n2253 VSS.t667 149.249
R1948 VSS.n2252 VSS.t523 149.249
R1949 VSS.n2251 VSS.t690 149.249
R1950 VSS.n2250 VSS.t519 149.249
R1951 VSS.n2249 VSS.t525 149.249
R1952 VSS.n2248 VSS.t605 149.249
R1953 VSS.n2247 VSS.t520 149.249
R1954 VSS.n2246 VSS.t602 149.249
R1955 VSS.n2245 VSS.t608 149.249
R1956 VSS.n2244 VSS.t708 149.249
R1957 VSS.n2243 VSS.t604 149.249
R1958 VSS.n2242 VSS.t705 149.249
R1959 VSS.n2241 VSS.t681 149.249
R1960 VSS.n2239 VSS.t675 149.249
R1961 VSS.n2238 VSS.t643 149.249
R1962 VSS.n2237 VSS.t538 149.249
R1963 VSS.n2236 VSS.t663 149.249
R1964 VSS.n2235 VSS.t746 149.249
R1965 VSS.n2234 VSS.t627 149.249
R1966 VSS.n2233 VSS.t513 149.249
R1967 VSS.n2232 VSS.t648 149.249
R1968 VSS.n2231 VSS.t722 149.249
R1969 VSS.n2230 VSS.t599 149.249
R1970 VSS.n2229 VSS.t660 149.249
R1971 VSS.n2228 VSS.t624 149.249
R1972 VSS.n2227 VSS.t621 149.249
R1973 VSS.n2226 VSS.t574 149.249
R1974 VSS.n2225 VSS.t644 149.249
R1975 VSS.n2159 VSS.t682 149.249
R1976 VSS.n2158 VSS.t655 149.249
R1977 VSS.n2157 VSS.t732 149.249
R1978 VSS.n2156 VSS.t612 149.249
R1979 VSS.n2155 VSS.t669 149.249
R1980 VSS.n2154 VSS.t635 149.249
R1981 VSS.n2153 VSS.t632 149.249
R1982 VSS.n2152 VSS.t583 149.249
R1983 VSS.n2151 VSS.t651 149.249
R1984 VSS.n2150 VSS.t611 149.249
R1985 VSS.n2149 VSS.t607 149.249
R1986 VSS.n2148 VSS.t728 149.249
R1987 VSS.n2147 VSS.t630 149.249
R1988 VSS.n2146 VSS.t750 149.249
R1989 VSS.n2145 VSS.t580 149.249
R1990 VSS.n2143 VSS.t548 149.249
R1991 VSS.n2142 VSS.t763 149.249
R1992 VSS.n2141 VSS.t662 149.249
R1993 VSS.n2140 VSS.t537 149.249
R1994 VSS.n2139 VSS.t625 149.249
R1995 VSS.n2138 VSS.t745 149.249
R1996 VSS.n2137 VSS.t647 149.249
R1997 VSS.n2136 VSS.t512 149.249
R1998 VSS.n2135 VSS.t597 149.249
R1999 VSS.n2134 VSS.t721 149.249
R2000 VSS.n2133 VSS.t532 149.249
R2001 VSS.n2132 VSS.t743 149.249
R2002 VSS.n2131 VSS.t740 149.249
R2003 VSS.n2130 VSS.t697 149.249
R2004 VSS.n2129 VSS.t764 149.249
R2005 VSS.n2029 VSS.t699 149.249
R2006 VSS.n2028 VSS.t671 149.249
R2007 VSS.n2027 VSS.t754 149.249
R2008 VSS.n2026 VSS.t634 149.249
R2009 VSS.n2025 VSS.t685 149.249
R2010 VSS.n2024 VSS.t653 149.249
R2011 VSS.n2023 VSS.t650 149.249
R2012 VSS.n2022 VSS.t610 149.249
R2013 VSS.n2021 VSS.t666 149.249
R2014 VSS.n2020 VSS.t631 149.249
R2015 VSS.n2019 VSS.t629 149.249
R2016 VSS.n2018 VSS.t749 149.249
R2017 VSS.n2017 VSS.t649 149.249
R2018 VSS.n2016 VSS.t518 149.249
R2019 VSS.n2015 VSS.t603 149.249
R2020 VSS.n2013 VSS.t564 149.249
R2021 VSS.n2012 VSS.t527 149.249
R2022 VSS.n2011 VSS.t679 149.249
R2023 VSS.n2010 VSS.t555 149.249
R2024 VSS.n2009 VSS.t646 149.249
R2025 VSS.n2008 VSS.t511 149.249
R2026 VSS.n2007 VSS.t659 149.249
R2027 VSS.n2006 VSS.t533 149.249
R2028 VSS.n2005 VSS.t620 149.249
R2029 VSS.n2004 VSS.t741 149.249
R2030 VSS.n2003 VSS.t549 149.249
R2031 VSS.n2002 VSS.t509 149.249
R2032 VSS.n2001 VSS.t759 149.249
R2033 VSS.n2000 VSS.t717 149.249
R2034 VSS.n1999 VSS.t528 149.249
R2035 VSS.n1933 VSS.t515 149.249
R2036 VSS.n1932 VSS.t733 149.249
R2037 VSS.n1931 VSS.t562 149.249
R2038 VSS.n1930 VSS.t688 149.249
R2039 VSS.n1929 VSS.t753 149.249
R2040 VSS.n1928 VSS.t709 149.249
R2041 VSS.n1927 VSS.t706 149.249
R2042 VSS.n1926 VSS.t668 149.249
R2043 VSS.n1925 VSS.t727 149.249
R2044 VSS.n1924 VSS.t686 149.249
R2045 VSS.n1923 VSS.t684 149.249
R2046 VSS.n1922 VSS.t561 149.249
R2047 VSS.n1921 VSS.t701 149.249
R2048 VSS.n1920 VSS.t581 149.249
R2049 VSS.n1919 VSS.t665 149.249
R2050 VSS.n1917 VSS.t638 149.249
R2051 VSS.n1916 VSS.t589 149.249
R2052 VSS.n1915 VSS.t744 149.249
R2053 VSS.n1914 VSS.t626 149.249
R2054 VSS.n1913 VSS.t698 149.249
R2055 VSS.n1912 VSS.t576 149.249
R2056 VSS.n1911 VSS.t720 149.249
R2057 VSS.n1910 VSS.t598 149.249
R2058 VSS.n1909 VSS.t677 149.249
R2059 VSS.n1908 VSS.t553 149.249
R2060 VSS.n1907 VSS.t619 149.249
R2061 VSS.n1906 VSS.t572 149.249
R2062 VSS.n1905 VSS.t568 149.249
R2063 VSS.n1904 VSS.t531 149.249
R2064 VSS.n1903 VSS.t591 149.249
R2065 VSS.n779 VSS.t617 149.249
R2066 VSS.n778 VSS.t579 149.249
R2067 VSS.n777 VSS.t664 149.249
R2068 VSS.n776 VSS.t540 149.249
R2069 VSS.n775 VSS.t601 149.249
R2070 VSS.n774 VSS.t559 149.249
R2071 VSS.n773 VSS.t557 149.249
R2072 VSS.n772 VSS.t514 149.249
R2073 VSS.n771 VSS.t577 149.249
R2074 VSS.n770 VSS.t536 149.249
R2075 VSS.n769 VSS.t535 149.249
R2076 VSS.n768 VSS.t661 149.249
R2077 VSS.n767 VSS.t554 149.249
R2078 VSS.n766 VSS.t678 149.249
R2079 VSS.n765 VSS.t510 149.249
R2080 VSS.n763 VSS.t640 149.249
R2081 VSS.n762 VSS.t593 149.249
R2082 VSS.n761 VSS.t747 149.249
R2083 VSS.n760 VSS.t628 149.249
R2084 VSS.n759 VSS.t700 149.249
R2085 VSS.n758 VSS.t578 149.249
R2086 VSS.n757 VSS.t723 149.249
R2087 VSS.n756 VSS.t600 149.249
R2088 VSS.n755 VSS.t680 149.249
R2089 VSS.n754 VSS.t556 149.249
R2090 VSS.n753 VSS.t622 149.249
R2091 VSS.n752 VSS.t575 149.249
R2092 VSS.n751 VSS.t571 149.249
R2093 VSS.n750 VSS.t534 149.249
R2094 VSS.n749 VSS.t594 149.249
R2095 VSS.n683 VSS.t539 149.249
R2096 VSS.n682 VSS.t758 149.249
R2097 VSS.n681 VSS.t584 149.249
R2098 VSS.n680 VSS.t710 149.249
R2099 VSS.n679 VSS.t522 149.249
R2100 VSS.n678 VSS.t731 149.249
R2101 VSS.n677 VSS.t730 149.249
R2102 VSS.n676 VSS.t687 149.249
R2103 VSS.n675 VSS.t752 149.249
R2104 VSS.n674 VSS.t707 149.249
R2105 VSS.n673 VSS.t704 149.249
R2106 VSS.n672 VSS.t582 149.249
R2107 VSS.n671 VSS.t726 149.249
R2108 VSS.n670 VSS.t606 149.249
R2109 VSS.n669 VSS.t683 149.249
R2110 VSS.n667 VSS.t558 149.249
R2111 VSS.n666 VSS.t516 149.249
R2112 VSS.n665 VSS.t670 149.249
R2113 VSS.n664 VSS.t545 149.249
R2114 VSS.n663 VSS.t633 149.249
R2115 VSS.n662 VSS.t755 149.249
R2116 VSS.n661 VSS.t652 149.249
R2117 VSS.n660 VSS.t521 149.249
R2118 VSS.n659 VSS.t609 149.249
R2119 VSS.n658 VSS.t729 149.249
R2120 VSS.n657 VSS.t543 149.249
R2121 VSS.n656 VSS.t751 149.249
R2122 VSS.n655 VSS.t748 149.249
R2123 VSS.n654 VSS.t703 149.249
R2124 VSS.n653 VSS.t517 149.249
R2125 VSS.n570 VSS.t524 149.249
R2126 VSS.n569 VSS.t742 149.249
R2127 VSS.n568 VSS.t570 149.249
R2128 VSS.n567 VSS.t695 149.249
R2129 VSS.n566 VSS.t761 149.249
R2130 VSS.n565 VSS.t718 149.249
R2131 VSS.n564 VSS.t715 149.249
R2132 VSS.n563 VSS.t676 149.249
R2133 VSS.n562 VSS.t736 149.249
R2134 VSS.n561 VSS.t694 149.249
R2135 VSS.n560 VSS.t692 149.249
R2136 VSS.n559 VSS.t565 149.249
R2137 VSS.n558 VSS.t712 149.249
R2138 VSS.n557 VSS.t585 149.249
R2139 VSS.n556 VSS.t673 149.249
R2140 VSS.n554 VSS.t544 149.249
R2141 VSS.n553 VSS.t756 149.249
R2142 VSS.n552 VSS.t657 149.249
R2143 VSS.n551 VSS.t529 149.249
R2144 VSS.n550 VSS.t616 149.249
R2145 VSS.n549 VSS.t737 149.249
R2146 VSS.n548 VSS.t639 149.249
R2147 VSS.n547 VSS.t760 149.249
R2148 VSS.n546 VSS.t588 149.249
R2149 VSS.n545 VSS.t714 149.249
R2150 VSS.n544 VSS.t526 149.249
R2151 VSS.n543 VSS.t735 149.249
R2152 VSS.n542 VSS.t734 149.249
R2153 VSS.n541 VSS.t691 149.249
R2154 VSS.n540 VSS.t757 149.249
R2155 VSS.n474 VSS.t654 149.249
R2156 VSS.n473 VSS.t623 149.249
R2157 VSS.n472 VSS.t696 149.249
R2158 VSS.n471 VSS.t573 149.249
R2159 VSS.n470 VSS.t642 149.249
R2160 VSS.n469 VSS.t595 149.249
R2161 VSS.n468 VSS.t592 149.249
R2162 VSS.n467 VSS.t551 149.249
R2163 VSS.n466 VSS.t615 149.249
R2164 VSS.n465 VSS.t569 149.249
R2165 VSS.n464 VSS.t567 149.249
R2166 VSS.n463 VSS.t693 149.249
R2167 VSS.n462 VSS.t587 149.249
R2168 VSS.n461 VSS.t713 149.249
R2169 VSS.n460 VSS.t547 149.249
R2170 VSS.n458 VSS.t672 149.249
R2171 VSS.n457 VSS.t636 149.249
R2172 VSS.n456 VSS.t530 149.249
R2173 VSS.n455 VSS.t658 149.249
R2174 VSS.n454 VSS.t739 149.249
R2175 VSS.n453 VSS.t618 149.249
R2176 VSS.n452 VSS.t762 149.249
R2177 VSS.n451 VSS.t641 149.249
R2178 VSS.n450 VSS.t716 149.249
R2179 VSS.n449 VSS.t590 149.249
R2180 VSS.n448 VSS.t656 149.249
R2181 VSS.n447 VSS.t614 149.249
R2182 VSS.n446 VSS.t613 149.249
R2183 VSS.n445 VSS.t566 149.249
R2184 VSS.n444 VSS.t637 149.249
R2185 VSS.n138 VSS.n137 145.921
R2186 VSS.n129 VSS.n128 145.921
R2187 VSS.n120 VSS.n119 145.921
R2188 VSS.n111 VSS.n110 145.921
R2189 VSS.n102 VSS.n101 145.921
R2190 VSS.n93 VSS.n92 145.921
R2191 VSS.n84 VSS.n83 145.921
R2192 VSS.n75 VSS.n74 145.921
R2193 VSS.n66 VSS.n65 145.921
R2194 VSS.n57 VSS.n56 145.921
R2195 VSS.n48 VSS.n47 145.921
R2196 VSS.n39 VSS.n38 145.921
R2197 VSS.n30 VSS.n29 145.921
R2198 VSS.n21 VSS.n20 145.921
R2199 VSS.n12 VSS.n11 145.921
R2200 VSS.n3 VSS.n2 145.921
R2201 VSS.n572 VSS.t2172 135.357
R2202 VSS.n1643 VSS.t1221 135.357
R2203 VSS.n575 VSS.t2415 135.357
R2204 VSS.n1112 VSS.t1285 135.357
R2205 VSS.n617 VSS.t2012 135.357
R2206 VSS.n1609 VSS.t486 135.357
R2207 VSS.n2092 VSS.t1688 135.357
R2208 VSS.n1080 VSS.t1548 135.357
R2209 VSS.n614 VSS.t1572 135.357
R2210 VSS.n1606 VSS.t2184 135.357
R2211 VSS.n2088 VSS.t2155 135.357
R2212 VSS.n1077 VSS.t1380 135.357
R2213 VSS.n611 VSS.t1375 135.357
R2214 VSS.n1603 VSS.t2519 135.357
R2215 VSS.n2084 VSS.t1743 135.357
R2216 VSS.n1074 VSS.t1853 135.357
R2217 VSS.n608 VSS.t1862 135.357
R2218 VSS.n1600 VSS.t2035 135.357
R2219 VSS.n2080 VSS.t2236 135.357
R2220 VSS.n1071 VSS.t1138 135.357
R2221 VSS.n605 VSS.t1104 135.357
R2222 VSS.n1597 VSS.t112 135.357
R2223 VSS.n2076 VSS.t2509 135.357
R2224 VSS.n1068 VSS.t995 135.357
R2225 VSS.n602 VSS.t1324 135.357
R2226 VSS.n1594 VSS.t2526 135.357
R2227 VSS.n2072 VSS.t1898 135.357
R2228 VSS.n1065 VSS.t818 135.357
R2229 VSS.n599 VSS.t899 135.357
R2230 VSS.n1591 VSS.t1435 135.357
R2231 VSS.n2068 VSS.t2139 135.357
R2232 VSS.n1062 VSS.t2292 135.357
R2233 VSS.n596 VSS.t2326 135.357
R2234 VSS.n1588 VSS.t2064 135.357
R2235 VSS.n2064 VSS.t811 135.357
R2236 VSS.n1059 VSS.t930 135.357
R2237 VSS.n593 VSS.t2422 135.357
R2238 VSS.n1585 VSS.t2107 135.357
R2239 VSS.n2060 VSS.t1603 135.357
R2240 VSS.n1056 VSS.t979 135.357
R2241 VSS.n590 VSS.t1055 135.357
R2242 VSS.n1582 VSS.t2372 135.357
R2243 VSS.n2056 VSS.t2374 135.357
R2244 VSS.n1053 VSS.t1631 135.357
R2245 VSS.n587 VSS.t2071 135.357
R2246 VSS.n1579 VSS.t1289 135.357
R2247 VSS.n2052 VSS.t400 135.357
R2248 VSS.n1050 VSS.t892 135.357
R2249 VSS.n584 VSS.t1112 135.357
R2250 VSS.n1576 VSS.t1737 135.357
R2251 VSS.n2048 VSS.t2191 135.357
R2252 VSS.n1047 VSS.t2242 135.357
R2253 VSS.n581 VSS.t1092 135.357
R2254 VSS.n1573 VSS.t880 135.357
R2255 VSS.n2044 VSS.t1994 135.357
R2256 VSS.n1044 VSS.t2027 135.357
R2257 VSS.n578 VSS.t1128 135.357
R2258 VSS.n1570 VSS.t967 135.357
R2259 VSS.n2040 VSS.t41 135.357
R2260 VSS.n1041 VSS.t1479 135.357
R2261 VSS.n1037 VSS.t769 135.357
R2262 VSS.n2036 VSS.t1678 135.357
R2263 VSS.n1567 VSS.t849 135.357
R2264 VSS.n2032 VSS.t2264 135.357
R2265 VSS.n411 VSS.t938 134.171
R2266 VSS.n410 VSS.t908 134.171
R2267 VSS.n407 VSS.t1694 134.171
R2268 VSS.n406 VSS.t2513 134.171
R2269 VSS.n403 VSS.t1999 134.171
R2270 VSS.n402 VSS.t802 134.171
R2271 VSS.n399 VSS.t1643 134.171
R2272 VSS.n398 VSS.t1784 134.171
R2273 VSS.n395 VSS.t1732 134.171
R2274 VSS.n394 VSS.t1174 134.171
R2275 VSS.n391 VSS.t446 134.171
R2276 VSS.n390 VSS.t2505 134.171
R2277 VSS.n387 VSS.t950 134.171
R2278 VSS.n386 VSS.t847 134.171
R2279 VSS.n383 VSS.t1814 134.171
R2280 VSS.n382 VSS.t973 134.171
R2281 VSS.n379 VSS.t1937 134.171
R2282 VSS.n378 VSS.t1248 134.171
R2283 VSS.n375 VSS.t2018 134.171
R2284 VSS.n374 VSS.t1764 134.171
R2285 VSS.n371 VSS.t1700 134.171
R2286 VSS.n370 VSS.t864 134.171
R2287 VSS.n367 VSS.t2116 134.171
R2288 VSS.n366 VSS.t2069 134.171
R2289 VSS.n363 VSS.t1353 134.171
R2290 VSS.n362 VSS.t1503 134.171
R2291 VSS.n359 VSS.t396 134.171
R2292 VSS.n358 VSS.t406 134.171
R2293 VSS.n355 VSS.t1281 134.171
R2294 VSS.n354 VSS.t1011 134.171
R2295 VSS.n351 VSS.t2356 134.171
R2296 VSS.n350 VSS.t2361 134.171
R2297 VSS.n2334 VSS.t134 125.574
R2298 VSS.n2331 VSS.t118 125.574
R2299 VSS.n2328 VSS.t132 125.574
R2300 VSS.n2325 VSS.t142 125.574
R2301 VSS.n2322 VSS.t148 125.574
R2302 VSS.n2319 VSS.t136 125.574
R2303 VSS.n2316 VSS.t122 125.574
R2304 VSS.n2313 VSS.t138 125.574
R2305 VSS.n2310 VSS.t120 125.574
R2306 VSS.n2307 VSS.t124 125.574
R2307 VSS.n2304 VSS.t140 125.574
R2308 VSS.n2301 VSS.t128 125.574
R2309 VSS.n2298 VSS.t126 125.574
R2310 VSS.n2295 VSS.t146 125.574
R2311 VSS.n2292 VSS.t130 125.574
R2312 VSS.n2289 VSS.t144 125.574
R2313 VSS.n2091 VSS.t233 89.332
R2314 VSS.n2087 VSS.t254 89.332
R2315 VSS.n2083 VSS.t151 89.332
R2316 VSS.n2079 VSS.t48 89.332
R2317 VSS.n2075 VSS.t260 89.332
R2318 VSS.n2071 VSS.t106 89.332
R2319 VSS.n2067 VSS.t0 89.332
R2320 VSS.n2063 VSS.t157 89.332
R2321 VSS.n2059 VSS.t39 89.332
R2322 VSS.n2055 VSS.t258 89.332
R2323 VSS.n2051 VSS.t238 89.332
R2324 VSS.n2047 VSS.t259 89.332
R2325 VSS.n2043 VSS.t255 89.332
R2326 VSS.n2039 VSS.t62 89.332
R2327 VSS.n2035 VSS.t257 89.332
R2328 VSS.n138 VSS.t95 76.337
R2329 VSS.n129 VSS.t1020 76.337
R2330 VSS.n120 VSS.t2434 76.337
R2331 VSS.n111 VSS.t1923 76.337
R2332 VSS.n102 VSS.t1574 76.337
R2333 VSS.n93 VSS.t2454 76.337
R2334 VSS.n84 VSS.t1082 76.337
R2335 VSS.n75 VSS.t98 76.337
R2336 VSS.n66 VSS.t780 76.337
R2337 VSS.n57 VSS.t1208 76.337
R2338 VSS.n48 VSS.t1154 76.337
R2339 VSS.n39 VSS.t983 76.337
R2340 VSS.n30 VSS.t2130 76.337
R2341 VSS.n21 VSS.t2313 76.337
R2342 VSS.n12 VSS.t2096 76.337
R2343 VSS.n3 VSS.t1395 76.337
R2344 VSS.t34 VSS.t70 68.097
R2345 VSS.t51 VSS.t26 68.097
R2346 VSS.t35 VSS.t11 68.097
R2347 VSS.t53 VSS.t8 68.097
R2348 VSS.t52 VSS.t7 68.097
R2349 VSS.t4 VSS.t24 68.097
R2350 VSS.t33 VSS.t9 68.097
R2351 VSS.t32 VSS.t18 68.097
R2352 VSS.t5 VSS.t25 68.097
R2353 VSS.t37 VSS.t29 68.097
R2354 VSS.t43 VSS.t75 68.097
R2355 VSS.t31 VSS.t72 68.097
R2356 VSS.t86 VSS.t23 68.097
R2357 VSS.t36 VSS.t15 68.097
R2358 VSS.t42 VSS.t27 68.097
R2359 VSS.t38 VSS.t21 68.097
R2360 VSS.t233 VSS.t68 65.168
R2361 VSS.t254 VSS.t74 65.168
R2362 VSS.t151 VSS.t71 65.168
R2363 VSS.t48 VSS.t20 65.168
R2364 VSS.t260 VSS.t14 65.168
R2365 VSS.t106 VSS.t17 65.168
R2366 VSS.t0 VSS.t54 65.168
R2367 VSS.t157 VSS.t19 65.168
R2368 VSS.t39 VSS.t12 65.168
R2369 VSS.t258 VSS.t69 65.168
R2370 VSS.t238 VSS.t28 65.168
R2371 VSS.t259 VSS.t73 65.168
R2372 VSS.t255 VSS.t22 65.168
R2373 VSS.t62 VSS.t16 65.168
R2374 VSS.t257 VSS.t13 65.168
R2375 VSS.t256 VSS.t10 65.168
R2376 VSS.n139 VSS.n138 63.013
R2377 VSS.n130 VSS.n129 63.013
R2378 VSS.n121 VSS.n120 63.013
R2379 VSS.n112 VSS.n111 63.013
R2380 VSS.n103 VSS.n102 63.013
R2381 VSS.n94 VSS.n93 63.013
R2382 VSS.n85 VSS.n84 63.013
R2383 VSS.n76 VSS.n75 63.013
R2384 VSS.n67 VSS.n66 63.013
R2385 VSS.n58 VSS.n57 63.013
R2386 VSS.n49 VSS.n48 63.013
R2387 VSS.n40 VSS.n39 63.013
R2388 VSS.n31 VSS.n30 63.013
R2389 VSS.n22 VSS.n21 63.013
R2390 VSS.n13 VSS.n12 63.013
R2391 VSS.n4 VSS.n3 63.013
R2392 VSS.n412 VSS.t1244 56.362
R2393 VSS.n408 VSS.t2524 56.362
R2394 VSS.n404 VSS.t1760 56.362
R2395 VSS.n400 VSS.t1423 56.362
R2396 VSS.n396 VSS.t1283 56.362
R2397 VSS.n392 VSS.t1235 56.362
R2398 VSS.n388 VSS.t1615 56.362
R2399 VSS.n384 VSS.t2016 56.362
R2400 VSS.n380 VSS.t1223 56.362
R2401 VSS.n376 VSS.t2103 56.362
R2402 VSS.n372 VSS.t1369 56.362
R2403 VSS.n368 VSS.t993 56.362
R2404 VSS.n364 VSS.t1691 56.362
R2405 VSS.n360 VSS.t1486 56.362
R2406 VSS.n356 VSS.t1714 56.362
R2407 VSS.n352 VSS.t1367 56.362
R2408 VSS.n350 VSS.t2402 55.057
R2409 VSS.n409 VSS.t910 53.505
R2410 VSS.n405 VSS.t2516 53.505
R2411 VSS.n401 VSS.t2275 53.505
R2412 VSS.n397 VSS.t957 53.505
R2413 VSS.n393 VSS.t1172 53.505
R2414 VSS.n389 VSS.t2507 53.505
R2415 VSS.n385 VSS.t845 53.505
R2416 VSS.n381 VSS.t1537 53.505
R2417 VSS.n377 VSS.t1246 53.505
R2418 VSS.n373 VSS.t1762 53.505
R2419 VSS.n369 VSS.t866 53.505
R2420 VSS.n365 VSS.t2067 53.505
R2421 VSS.n361 VSS.t1501 53.505
R2422 VSS.n357 VSS.t403 53.505
R2423 VSS.n353 VSS.t1009 53.505
R2424 VSS.t332 VSS.t2225 44.494
R2425 VSS.t366 VSS.t2234 44.494
R2426 VSS.t341 VSS.t2227 44.494
R2427 VSS.t365 VSS.t2233 44.494
R2428 VSS.t363 VSS.t2232 44.494
R2429 VSS.t279 VSS.t2220 44.494
R2430 VSS.t297 VSS.t2223 44.494
R2431 VSS.t347 VSS.t2230 44.494
R2432 VSS.t296 VSS.t2222 44.494
R2433 VSS.t346 VSS.t2229 44.494
R2434 VSS.t291 VSS.t2221 44.494
R2435 VSS.t342 VSS.t2228 44.494
R2436 VSS.t357 VSS.t2231 44.494
R2437 VSS.t361 VSS.t1922 44.494
R2438 VSS.t368 VSS.t2433 44.494
R2439 VSS.t326 VSS.t1019 44.494
R2440 VSS.t277 VSS.t91 44.494
R2441 VSS.t308 VSS.t1984 44.494
R2442 VSS.t348 VSS.t832 44.494
R2443 VSS.t315 VSS.t825 44.494
R2444 VSS.t345 VSS.t831 44.494
R2445 VSS.t340 VSS.t830 44.494
R2446 VSS.t370 VSS.t1979 44.494
R2447 VSS.t276 VSS.t1982 44.494
R2448 VSS.t322 VSS.t828 44.494
R2449 VSS.t275 VSS.t1981 44.494
R2450 VSS.t320 VSS.t827 44.494
R2451 VSS.t271 VSS.t1980 44.494
R2452 VSS.t318 VSS.t826 44.494
R2453 VSS.t331 VSS.t829 44.494
R2454 VSS.t338 VSS.t1924 44.494
R2455 VSS.t350 VSS.t2436 44.494
R2456 VSS.t302 VSS.t1021 44.494
R2457 VSS.t262 VSS.t2 44.494
R2458 VSS.n2126 VSS.n2034 43.368
R2459 VSS.n2124 VSS.n2038 43.368
R2460 VSS.n2122 VSS.n2042 43.368
R2461 VSS.n2120 VSS.n2046 43.368
R2462 VSS.n2118 VSS.n2050 43.368
R2463 VSS.n2116 VSS.n2054 43.368
R2464 VSS.n2114 VSS.n2058 43.368
R2465 VSS.n2112 VSS.n2062 43.368
R2466 VSS.n2110 VSS.n2066 43.368
R2467 VSS.n2108 VSS.n2070 43.368
R2468 VSS.n2106 VSS.n2074 43.368
R2469 VSS.n2104 VSS.n2078 43.368
R2470 VSS.n2102 VSS.n2082 43.368
R2471 VSS.n2100 VSS.n2086 43.368
R2472 VSS.n2098 VSS.n2090 43.368
R2473 VSS.t266 VSS.t1394 42.022
R2474 VSS.t294 VSS.t2095 42.022
R2475 VSS.t304 VSS.t2312 42.022
R2476 VSS.t313 VSS.t2129 42.022
R2477 VSS.t323 VSS.t982 42.022
R2478 VSS.t309 VSS.t1153 42.022
R2479 VSS.t269 VSS.t1207 42.022
R2480 VSS.t306 VSS.t779 42.022
R2481 VSS.t359 VSS.t97 42.022
R2482 VSS.t264 VSS.t495 42.022
R2483 VSS.t354 VSS.t2453 42.022
R2484 VSS.t316 VSS.t1573 42.022
R2485 VSS.t325 VSS.t2224 42.022
R2486 VSS.t268 VSS.t2219 42.022
R2487 VSS.t336 VSS.t2226 42.022
R2488 VSS.t376 VSS.t1396 42.022
R2489 VSS.t273 VSS.t2098 42.022
R2490 VSS.t281 VSS.t2315 42.022
R2491 VSS.t289 VSS.t2132 42.022
R2492 VSS.t298 VSS.t984 42.022
R2493 VSS.t286 VSS.t1156 42.022
R2494 VSS.t378 VSS.t1209 42.022
R2495 VSS.t284 VSS.t782 42.022
R2496 VSS.t333 VSS.t99 42.022
R2497 VSS.t372 VSS.t1064 42.022
R2498 VSS.t329 VSS.t2456 42.022
R2499 VSS.t292 VSS.t1575 42.022
R2500 VSS.t301 VSS.t1983 42.022
R2501 VSS.t364 VSS.t1978 42.022
R2502 VSS.t312 VSS.t824 42.022
R2503 VSS.n650 VSS.n574 41.109
R2504 VSS.n648 VSS.n577 41.109
R2505 VSS.n646 VSS.n580 41.109
R2506 VSS.n644 VSS.n583 41.109
R2507 VSS.n642 VSS.n586 41.109
R2508 VSS.n640 VSS.n589 41.109
R2509 VSS.n638 VSS.n592 41.109
R2510 VSS.n636 VSS.n595 41.109
R2511 VSS.n634 VSS.n598 41.109
R2512 VSS.n632 VSS.n601 41.109
R2513 VSS.n630 VSS.n604 41.109
R2514 VSS.n628 VSS.n607 41.109
R2515 VSS.n626 VSS.n610 41.109
R2516 VSS.n624 VSS.n613 41.109
R2517 VSS.n622 VSS.n616 41.109
R2518 VSS.n305 VSS.t301 39.55
R2519 VSS.n314 VSS.t364 39.55
R2520 VSS.n323 VSS.t312 39.55
R2521 VSS.n189 VSS.t308 37.078
R2522 VSS.n197 VSS.t348 37.078
R2523 VSS.n206 VSS.t315 37.078
R2524 VSS.n215 VSS.t345 37.078
R2525 VSS.n224 VSS.t340 37.078
R2526 VSS.n233 VSS.t370 37.078
R2527 VSS.n242 VSS.t276 37.078
R2528 VSS.n251 VSS.t322 37.078
R2529 VSS.n260 VSS.t275 37.078
R2530 VSS.n269 VSS.t320 37.078
R2531 VSS.n278 VSS.t271 37.078
R2532 VSS.n287 VSS.t318 37.078
R2533 VSS.n296 VSS.t331 37.078
R2534 VSS.n2096 VSS.n2094 32.376
R2535 VSS.n2095 VSS.t256 31.486
R2536 VSS.n620 VSS.n619 30.117
R2537 VSS.n1642 VSS.n1566 29.815
R2538 VSS.n1640 VSS.n1569 29.815
R2539 VSS.n1638 VSS.n1572 29.815
R2540 VSS.n1636 VSS.n1575 29.815
R2541 VSS.n1634 VSS.n1578 29.815
R2542 VSS.n1632 VSS.n1581 29.815
R2543 VSS.n1630 VSS.n1584 29.815
R2544 VSS.n1628 VSS.n1587 29.815
R2545 VSS.n1626 VSS.n1590 29.815
R2546 VSS.n1624 VSS.n1593 29.815
R2547 VSS.n1622 VSS.n1596 29.815
R2548 VSS.n1620 VSS.n1599 29.815
R2549 VSS.n1618 VSS.n1602 29.815
R2550 VSS.n1616 VSS.n1605 29.815
R2551 VSS.n1614 VSS.n1608 29.815
R2552 VSS.n1115 VSS.n1039 29.062
R2553 VSS.n1111 VSS.n1040 29.062
R2554 VSS.n1109 VSS.n1043 29.062
R2555 VSS.n1107 VSS.n1046 29.062
R2556 VSS.n1105 VSS.n1049 29.062
R2557 VSS.n1103 VSS.n1052 29.062
R2558 VSS.n1101 VSS.n1055 29.062
R2559 VSS.n1099 VSS.n1058 29.062
R2560 VSS.n1097 VSS.n1061 29.062
R2561 VSS.n1095 VSS.n1064 29.062
R2562 VSS.n1093 VSS.n1067 29.062
R2563 VSS.n1091 VSS.n1070 29.062
R2564 VSS.n1089 VSS.n1073 29.062
R2565 VSS.n1087 VSS.n1076 29.062
R2566 VSS.n1085 VSS.n1079 29.062
R2567 VSS.n415 VSS.n413 27.69
R2568 VSS.n573 VSS.n572 27.367
R2569 VSS.n576 VSS.n575 27.367
R2570 VSS.n618 VSS.n617 27.367
R2571 VSS.n1610 VSS.n1609 27.367
R2572 VSS.n2093 VSS.n2092 27.367
R2573 VSS.n1081 VSS.n1080 27.367
R2574 VSS.n615 VSS.n614 27.367
R2575 VSS.n1607 VSS.n1606 27.367
R2576 VSS.n2089 VSS.n2088 27.367
R2577 VSS.n1078 VSS.n1077 27.367
R2578 VSS.n612 VSS.n611 27.367
R2579 VSS.n1604 VSS.n1603 27.367
R2580 VSS.n2085 VSS.n2084 27.367
R2581 VSS.n1075 VSS.n1074 27.367
R2582 VSS.n609 VSS.n608 27.367
R2583 VSS.n1601 VSS.n1600 27.367
R2584 VSS.n2081 VSS.n2080 27.367
R2585 VSS.n1072 VSS.n1071 27.367
R2586 VSS.n606 VSS.n605 27.367
R2587 VSS.n1598 VSS.n1597 27.367
R2588 VSS.n2077 VSS.n2076 27.367
R2589 VSS.n1069 VSS.n1068 27.367
R2590 VSS.n603 VSS.n602 27.367
R2591 VSS.n1595 VSS.n1594 27.367
R2592 VSS.n2073 VSS.n2072 27.367
R2593 VSS.n1066 VSS.n1065 27.367
R2594 VSS.n600 VSS.n599 27.367
R2595 VSS.n1592 VSS.n1591 27.367
R2596 VSS.n2069 VSS.n2068 27.367
R2597 VSS.n1063 VSS.n1062 27.367
R2598 VSS.n597 VSS.n596 27.367
R2599 VSS.n1589 VSS.n1588 27.367
R2600 VSS.n2065 VSS.n2064 27.367
R2601 VSS.n1060 VSS.n1059 27.367
R2602 VSS.n594 VSS.n593 27.367
R2603 VSS.n1586 VSS.n1585 27.367
R2604 VSS.n2061 VSS.n2060 27.367
R2605 VSS.n1057 VSS.n1056 27.367
R2606 VSS.n591 VSS.n590 27.367
R2607 VSS.n1583 VSS.n1582 27.367
R2608 VSS.n2057 VSS.n2056 27.367
R2609 VSS.n1054 VSS.n1053 27.367
R2610 VSS.n588 VSS.n587 27.367
R2611 VSS.n1580 VSS.n1579 27.367
R2612 VSS.n2053 VSS.n2052 27.367
R2613 VSS.n1051 VSS.n1050 27.367
R2614 VSS.n585 VSS.n584 27.367
R2615 VSS.n1577 VSS.n1576 27.367
R2616 VSS.n2049 VSS.n2048 27.367
R2617 VSS.n1048 VSS.n1047 27.367
R2618 VSS.n582 VSS.n581 27.367
R2619 VSS.n1574 VSS.n1573 27.367
R2620 VSS.n2045 VSS.n2044 27.367
R2621 VSS.n1045 VSS.n1044 27.367
R2622 VSS.n579 VSS.n578 27.367
R2623 VSS.n1571 VSS.n1570 27.367
R2624 VSS.n2041 VSS.n2040 27.367
R2625 VSS.n1042 VSS.n1041 27.367
R2626 VSS.n1038 VSS.n1037 27.367
R2627 VSS.n1113 VSS.n1112 27.367
R2628 VSS.n2037 VSS.n2036 27.367
R2629 VSS.n1568 VSS.n1567 27.367
R2630 VSS.n1644 VSS.n1643 27.367
R2631 VSS.n2033 VSS.n2032 27.367
R2632 VSS.n2338 VSS.n334 27.194
R2633 VSS.n116 VSS.t325 27.191
R2634 VSS.n125 VSS.t268 27.191
R2635 VSS.n134 VSS.t336 27.191
R2636 VSS.n2178 VSS.n2177 25.944
R2637 VSS.n1952 VSS.n1951 25.944
R2638 VSS.n1856 VSS.n1855 25.944
R2639 VSS.n1792 VSS.n1791 25.944
R2640 VSS.n1728 VSS.n1727 25.944
R2641 VSS.n1664 VSS.n1663 25.944
R2642 VSS.n1519 VSS.n1518 25.944
R2643 VSS.n1455 VSS.n1454 25.944
R2644 VSS.n1391 VSS.n1390 25.944
R2645 VSS.n1327 VSS.n1326 25.944
R2646 VSS.n1263 VSS.n1262 25.944
R2647 VSS.n1199 VSS.n1198 25.944
R2648 VSS.n1135 VSS.n1134 25.944
R2649 VSS.n990 VSS.n989 25.944
R2650 VSS.n926 VSS.n925 25.944
R2651 VSS.n862 VSS.n861 25.944
R2652 VSS.n798 VSS.n797 25.944
R2653 VSS.n702 VSS.n701 25.944
R2654 VSS.n493 VSS.n492 25.944
R2655 VSS.n0 VSS.t332 24.719
R2656 VSS.n8 VSS.t366 24.719
R2657 VSS.n17 VSS.t341 24.719
R2658 VSS.n26 VSS.t365 24.719
R2659 VSS.n35 VSS.t363 24.719
R2660 VSS.n44 VSS.t279 24.719
R2661 VSS.n53 VSS.t297 24.719
R2662 VSS.n62 VSS.t347 24.719
R2663 VSS.n71 VSS.t296 24.719
R2664 VSS.n80 VSS.t346 24.719
R2665 VSS.n89 VSS.t291 24.719
R2666 VSS.n98 VSS.t342 24.719
R2667 VSS.n107 VSS.t357 24.719
R2668 VSS.n343 VSS.n342 24.468
R2669 VSS.n1 VSS.n0 24.372
R2670 VSS.n9 VSS.n8 24.372
R2671 VSS.n18 VSS.n17 24.372
R2672 VSS.n27 VSS.n26 24.372
R2673 VSS.n36 VSS.n35 24.372
R2674 VSS.n45 VSS.n44 24.372
R2675 VSS.n54 VSS.n53 24.372
R2676 VSS.n63 VSS.n62 24.372
R2677 VSS.n72 VSS.n71 24.372
R2678 VSS.n81 VSS.n80 24.372
R2679 VSS.n90 VSS.n89 24.372
R2680 VSS.n99 VSS.n98 24.372
R2681 VSS.n108 VSS.n107 24.372
R2682 VSS.n117 VSS.n116 24.372
R2683 VSS.n126 VSS.n125 24.372
R2684 VSS.n135 VSS.n134 24.372
R2685 VSS.n2291 VSS.n2290 22.959
R2686 VSS.n2294 VSS.n2293 22.959
R2687 VSS.n2297 VSS.n2296 22.959
R2688 VSS.n2300 VSS.n2299 22.959
R2689 VSS.n2303 VSS.n2302 22.959
R2690 VSS.n2306 VSS.n2305 22.959
R2691 VSS.n2309 VSS.n2308 22.959
R2692 VSS.n2312 VSS.n2311 22.959
R2693 VSS.n2315 VSS.n2314 22.959
R2694 VSS.n2318 VSS.n2317 22.959
R2695 VSS.n2321 VSS.n2320 22.959
R2696 VSS.n2324 VSS.n2323 22.959
R2697 VSS.n2327 VSS.n2326 22.959
R2698 VSS.n2330 VSS.n2329 22.959
R2699 VSS.n2333 VSS.n2332 22.959
R2700 VSS.n190 VSS.n189 22.885
R2701 VSS.n198 VSS.n197 22.885
R2702 VSS.n207 VSS.n206 22.885
R2703 VSS.n216 VSS.n215 22.885
R2704 VSS.n225 VSS.n224 22.885
R2705 VSS.n234 VSS.n233 22.885
R2706 VSS.n243 VSS.n242 22.885
R2707 VSS.n252 VSS.n251 22.885
R2708 VSS.n261 VSS.n260 22.885
R2709 VSS.n270 VSS.n269 22.885
R2710 VSS.n279 VSS.n278 22.885
R2711 VSS.n288 VSS.n287 22.885
R2712 VSS.n297 VSS.n296 22.885
R2713 VSS.n306 VSS.n305 22.885
R2714 VSS.n315 VSS.n314 22.885
R2715 VSS.n324 VSS.n323 22.885
R2716 VSS.n2222 VSS.n2221 22.72
R2717 VSS.n2219 VSS.n2218 22.72
R2718 VSS.n2216 VSS.n2215 22.72
R2719 VSS.n2213 VSS.n2212 22.72
R2720 VSS.n2210 VSS.n2209 22.72
R2721 VSS.n2207 VSS.n2206 22.72
R2722 VSS.n2204 VSS.n2203 22.72
R2723 VSS.n2201 VSS.n2200 22.72
R2724 VSS.n2198 VSS.n2197 22.72
R2725 VSS.n2195 VSS.n2194 22.72
R2726 VSS.n2192 VSS.n2191 22.72
R2727 VSS.n2189 VSS.n2188 22.72
R2728 VSS.n2186 VSS.n2185 22.72
R2729 VSS.n2183 VSS.n2182 22.72
R2730 VSS.n2180 VSS.n2179 22.72
R2731 VSS.n1996 VSS.n1995 22.72
R2732 VSS.n1993 VSS.n1992 22.72
R2733 VSS.n1990 VSS.n1989 22.72
R2734 VSS.n1987 VSS.n1986 22.72
R2735 VSS.n1984 VSS.n1983 22.72
R2736 VSS.n1981 VSS.n1980 22.72
R2737 VSS.n1978 VSS.n1977 22.72
R2738 VSS.n1975 VSS.n1974 22.72
R2739 VSS.n1972 VSS.n1971 22.72
R2740 VSS.n1969 VSS.n1968 22.72
R2741 VSS.n1966 VSS.n1965 22.72
R2742 VSS.n1963 VSS.n1962 22.72
R2743 VSS.n1960 VSS.n1959 22.72
R2744 VSS.n1957 VSS.n1956 22.72
R2745 VSS.n1954 VSS.n1953 22.72
R2746 VSS.n1900 VSS.n1899 22.72
R2747 VSS.n1897 VSS.n1896 22.72
R2748 VSS.n1894 VSS.n1893 22.72
R2749 VSS.n1891 VSS.n1890 22.72
R2750 VSS.n1888 VSS.n1887 22.72
R2751 VSS.n1885 VSS.n1884 22.72
R2752 VSS.n1882 VSS.n1881 22.72
R2753 VSS.n1879 VSS.n1878 22.72
R2754 VSS.n1876 VSS.n1875 22.72
R2755 VSS.n1873 VSS.n1872 22.72
R2756 VSS.n1870 VSS.n1869 22.72
R2757 VSS.n1867 VSS.n1866 22.72
R2758 VSS.n1864 VSS.n1863 22.72
R2759 VSS.n1861 VSS.n1860 22.72
R2760 VSS.n1858 VSS.n1857 22.72
R2761 VSS.n1836 VSS.n1835 22.72
R2762 VSS.n1833 VSS.n1832 22.72
R2763 VSS.n1830 VSS.n1829 22.72
R2764 VSS.n1827 VSS.n1826 22.72
R2765 VSS.n1824 VSS.n1823 22.72
R2766 VSS.n1821 VSS.n1820 22.72
R2767 VSS.n1818 VSS.n1817 22.72
R2768 VSS.n1815 VSS.n1814 22.72
R2769 VSS.n1812 VSS.n1811 22.72
R2770 VSS.n1809 VSS.n1808 22.72
R2771 VSS.n1806 VSS.n1805 22.72
R2772 VSS.n1803 VSS.n1802 22.72
R2773 VSS.n1800 VSS.n1799 22.72
R2774 VSS.n1797 VSS.n1796 22.72
R2775 VSS.n1794 VSS.n1793 22.72
R2776 VSS.n1772 VSS.n1771 22.72
R2777 VSS.n1769 VSS.n1768 22.72
R2778 VSS.n1766 VSS.n1765 22.72
R2779 VSS.n1763 VSS.n1762 22.72
R2780 VSS.n1760 VSS.n1759 22.72
R2781 VSS.n1757 VSS.n1756 22.72
R2782 VSS.n1754 VSS.n1753 22.72
R2783 VSS.n1751 VSS.n1750 22.72
R2784 VSS.n1748 VSS.n1747 22.72
R2785 VSS.n1745 VSS.n1744 22.72
R2786 VSS.n1742 VSS.n1741 22.72
R2787 VSS.n1739 VSS.n1738 22.72
R2788 VSS.n1736 VSS.n1735 22.72
R2789 VSS.n1733 VSS.n1732 22.72
R2790 VSS.n1730 VSS.n1729 22.72
R2791 VSS.n1708 VSS.n1707 22.72
R2792 VSS.n1705 VSS.n1704 22.72
R2793 VSS.n1702 VSS.n1701 22.72
R2794 VSS.n1699 VSS.n1698 22.72
R2795 VSS.n1696 VSS.n1695 22.72
R2796 VSS.n1693 VSS.n1692 22.72
R2797 VSS.n1690 VSS.n1689 22.72
R2798 VSS.n1687 VSS.n1686 22.72
R2799 VSS.n1684 VSS.n1683 22.72
R2800 VSS.n1681 VSS.n1680 22.72
R2801 VSS.n1678 VSS.n1677 22.72
R2802 VSS.n1675 VSS.n1674 22.72
R2803 VSS.n1672 VSS.n1671 22.72
R2804 VSS.n1669 VSS.n1668 22.72
R2805 VSS.n1666 VSS.n1665 22.72
R2806 VSS.n1563 VSS.n1562 22.72
R2807 VSS.n1560 VSS.n1559 22.72
R2808 VSS.n1557 VSS.n1556 22.72
R2809 VSS.n1554 VSS.n1553 22.72
R2810 VSS.n1551 VSS.n1550 22.72
R2811 VSS.n1548 VSS.n1547 22.72
R2812 VSS.n1545 VSS.n1544 22.72
R2813 VSS.n1542 VSS.n1541 22.72
R2814 VSS.n1539 VSS.n1538 22.72
R2815 VSS.n1536 VSS.n1535 22.72
R2816 VSS.n1533 VSS.n1532 22.72
R2817 VSS.n1530 VSS.n1529 22.72
R2818 VSS.n1527 VSS.n1526 22.72
R2819 VSS.n1524 VSS.n1523 22.72
R2820 VSS.n1521 VSS.n1520 22.72
R2821 VSS.n1499 VSS.n1498 22.72
R2822 VSS.n1496 VSS.n1495 22.72
R2823 VSS.n1493 VSS.n1492 22.72
R2824 VSS.n1490 VSS.n1489 22.72
R2825 VSS.n1487 VSS.n1486 22.72
R2826 VSS.n1484 VSS.n1483 22.72
R2827 VSS.n1481 VSS.n1480 22.72
R2828 VSS.n1478 VSS.n1477 22.72
R2829 VSS.n1475 VSS.n1474 22.72
R2830 VSS.n1472 VSS.n1471 22.72
R2831 VSS.n1469 VSS.n1468 22.72
R2832 VSS.n1466 VSS.n1465 22.72
R2833 VSS.n1463 VSS.n1462 22.72
R2834 VSS.n1460 VSS.n1459 22.72
R2835 VSS.n1457 VSS.n1456 22.72
R2836 VSS.n1435 VSS.n1434 22.72
R2837 VSS.n1432 VSS.n1431 22.72
R2838 VSS.n1429 VSS.n1428 22.72
R2839 VSS.n1426 VSS.n1425 22.72
R2840 VSS.n1423 VSS.n1422 22.72
R2841 VSS.n1420 VSS.n1419 22.72
R2842 VSS.n1417 VSS.n1416 22.72
R2843 VSS.n1414 VSS.n1413 22.72
R2844 VSS.n1411 VSS.n1410 22.72
R2845 VSS.n1408 VSS.n1407 22.72
R2846 VSS.n1405 VSS.n1404 22.72
R2847 VSS.n1402 VSS.n1401 22.72
R2848 VSS.n1399 VSS.n1398 22.72
R2849 VSS.n1396 VSS.n1395 22.72
R2850 VSS.n1393 VSS.n1392 22.72
R2851 VSS.n1371 VSS.n1370 22.72
R2852 VSS.n1368 VSS.n1367 22.72
R2853 VSS.n1365 VSS.n1364 22.72
R2854 VSS.n1362 VSS.n1361 22.72
R2855 VSS.n1359 VSS.n1358 22.72
R2856 VSS.n1356 VSS.n1355 22.72
R2857 VSS.n1353 VSS.n1352 22.72
R2858 VSS.n1350 VSS.n1349 22.72
R2859 VSS.n1347 VSS.n1346 22.72
R2860 VSS.n1344 VSS.n1343 22.72
R2861 VSS.n1341 VSS.n1340 22.72
R2862 VSS.n1338 VSS.n1337 22.72
R2863 VSS.n1335 VSS.n1334 22.72
R2864 VSS.n1332 VSS.n1331 22.72
R2865 VSS.n1329 VSS.n1328 22.72
R2866 VSS.n1307 VSS.n1306 22.72
R2867 VSS.n1304 VSS.n1303 22.72
R2868 VSS.n1301 VSS.n1300 22.72
R2869 VSS.n1298 VSS.n1297 22.72
R2870 VSS.n1295 VSS.n1294 22.72
R2871 VSS.n1292 VSS.n1291 22.72
R2872 VSS.n1289 VSS.n1288 22.72
R2873 VSS.n1286 VSS.n1285 22.72
R2874 VSS.n1283 VSS.n1282 22.72
R2875 VSS.n1280 VSS.n1279 22.72
R2876 VSS.n1277 VSS.n1276 22.72
R2877 VSS.n1274 VSS.n1273 22.72
R2878 VSS.n1271 VSS.n1270 22.72
R2879 VSS.n1268 VSS.n1267 22.72
R2880 VSS.n1265 VSS.n1264 22.72
R2881 VSS.n1243 VSS.n1242 22.72
R2882 VSS.n1240 VSS.n1239 22.72
R2883 VSS.n1237 VSS.n1236 22.72
R2884 VSS.n1234 VSS.n1233 22.72
R2885 VSS.n1231 VSS.n1230 22.72
R2886 VSS.n1228 VSS.n1227 22.72
R2887 VSS.n1225 VSS.n1224 22.72
R2888 VSS.n1222 VSS.n1221 22.72
R2889 VSS.n1219 VSS.n1218 22.72
R2890 VSS.n1216 VSS.n1215 22.72
R2891 VSS.n1213 VSS.n1212 22.72
R2892 VSS.n1210 VSS.n1209 22.72
R2893 VSS.n1207 VSS.n1206 22.72
R2894 VSS.n1204 VSS.n1203 22.72
R2895 VSS.n1201 VSS.n1200 22.72
R2896 VSS.n1179 VSS.n1178 22.72
R2897 VSS.n1176 VSS.n1175 22.72
R2898 VSS.n1173 VSS.n1172 22.72
R2899 VSS.n1170 VSS.n1169 22.72
R2900 VSS.n1167 VSS.n1166 22.72
R2901 VSS.n1164 VSS.n1163 22.72
R2902 VSS.n1161 VSS.n1160 22.72
R2903 VSS.n1158 VSS.n1157 22.72
R2904 VSS.n1155 VSS.n1154 22.72
R2905 VSS.n1152 VSS.n1151 22.72
R2906 VSS.n1149 VSS.n1148 22.72
R2907 VSS.n1146 VSS.n1145 22.72
R2908 VSS.n1143 VSS.n1142 22.72
R2909 VSS.n1140 VSS.n1139 22.72
R2910 VSS.n1137 VSS.n1136 22.72
R2911 VSS.n1034 VSS.n1033 22.72
R2912 VSS.n1031 VSS.n1030 22.72
R2913 VSS.n1028 VSS.n1027 22.72
R2914 VSS.n1025 VSS.n1024 22.72
R2915 VSS.n1022 VSS.n1021 22.72
R2916 VSS.n1019 VSS.n1018 22.72
R2917 VSS.n1016 VSS.n1015 22.72
R2918 VSS.n1013 VSS.n1012 22.72
R2919 VSS.n1010 VSS.n1009 22.72
R2920 VSS.n1007 VSS.n1006 22.72
R2921 VSS.n1004 VSS.n1003 22.72
R2922 VSS.n1001 VSS.n1000 22.72
R2923 VSS.n998 VSS.n997 22.72
R2924 VSS.n995 VSS.n994 22.72
R2925 VSS.n992 VSS.n991 22.72
R2926 VSS.n970 VSS.n969 22.72
R2927 VSS.n967 VSS.n966 22.72
R2928 VSS.n964 VSS.n963 22.72
R2929 VSS.n961 VSS.n960 22.72
R2930 VSS.n958 VSS.n957 22.72
R2931 VSS.n955 VSS.n954 22.72
R2932 VSS.n952 VSS.n951 22.72
R2933 VSS.n949 VSS.n948 22.72
R2934 VSS.n946 VSS.n945 22.72
R2935 VSS.n943 VSS.n942 22.72
R2936 VSS.n940 VSS.n939 22.72
R2937 VSS.n937 VSS.n936 22.72
R2938 VSS.n934 VSS.n933 22.72
R2939 VSS.n931 VSS.n930 22.72
R2940 VSS.n928 VSS.n927 22.72
R2941 VSS.n906 VSS.n905 22.72
R2942 VSS.n903 VSS.n902 22.72
R2943 VSS.n900 VSS.n899 22.72
R2944 VSS.n897 VSS.n896 22.72
R2945 VSS.n894 VSS.n893 22.72
R2946 VSS.n891 VSS.n890 22.72
R2947 VSS.n888 VSS.n887 22.72
R2948 VSS.n885 VSS.n884 22.72
R2949 VSS.n882 VSS.n881 22.72
R2950 VSS.n879 VSS.n878 22.72
R2951 VSS.n876 VSS.n875 22.72
R2952 VSS.n873 VSS.n872 22.72
R2953 VSS.n870 VSS.n869 22.72
R2954 VSS.n867 VSS.n866 22.72
R2955 VSS.n864 VSS.n863 22.72
R2956 VSS.n842 VSS.n841 22.72
R2957 VSS.n839 VSS.n838 22.72
R2958 VSS.n836 VSS.n835 22.72
R2959 VSS.n833 VSS.n832 22.72
R2960 VSS.n830 VSS.n829 22.72
R2961 VSS.n827 VSS.n826 22.72
R2962 VSS.n824 VSS.n823 22.72
R2963 VSS.n821 VSS.n820 22.72
R2964 VSS.n818 VSS.n817 22.72
R2965 VSS.n815 VSS.n814 22.72
R2966 VSS.n812 VSS.n811 22.72
R2967 VSS.n809 VSS.n808 22.72
R2968 VSS.n806 VSS.n805 22.72
R2969 VSS.n803 VSS.n802 22.72
R2970 VSS.n800 VSS.n799 22.72
R2971 VSS.n746 VSS.n745 22.72
R2972 VSS.n743 VSS.n742 22.72
R2973 VSS.n740 VSS.n739 22.72
R2974 VSS.n737 VSS.n736 22.72
R2975 VSS.n734 VSS.n733 22.72
R2976 VSS.n731 VSS.n730 22.72
R2977 VSS.n728 VSS.n727 22.72
R2978 VSS.n725 VSS.n724 22.72
R2979 VSS.n722 VSS.n721 22.72
R2980 VSS.n719 VSS.n718 22.72
R2981 VSS.n716 VSS.n715 22.72
R2982 VSS.n713 VSS.n712 22.72
R2983 VSS.n710 VSS.n709 22.72
R2984 VSS.n707 VSS.n706 22.72
R2985 VSS.n704 VSS.n703 22.72
R2986 VSS.n537 VSS.n536 22.72
R2987 VSS.n534 VSS.n533 22.72
R2988 VSS.n531 VSS.n530 22.72
R2989 VSS.n528 VSS.n527 22.72
R2990 VSS.n525 VSS.n524 22.72
R2991 VSS.n522 VSS.n521 22.72
R2992 VSS.n519 VSS.n518 22.72
R2993 VSS.n516 VSS.n515 22.72
R2994 VSS.n513 VSS.n512 22.72
R2995 VSS.n510 VSS.n509 22.72
R2996 VSS.n507 VSS.n506 22.72
R2997 VSS.n504 VSS.n503 22.72
R2998 VSS.n501 VSS.n500 22.72
R2999 VSS.n498 VSS.n497 22.72
R3000 VSS.n495 VSS.n494 22.72
R3001 VSS.n443 VSS.n442 22.72
R3002 VSS.n441 VSS.n440 22.72
R3003 VSS.n439 VSS.n438 22.72
R3004 VSS.n437 VSS.n436 22.72
R3005 VSS.n435 VSS.n434 22.72
R3006 VSS.n433 VSS.n432 22.72
R3007 VSS.n431 VSS.n430 22.72
R3008 VSS.n429 VSS.n428 22.72
R3009 VSS.n427 VSS.n426 22.72
R3010 VSS.n425 VSS.n424 22.72
R3011 VSS.n423 VSS.n422 22.72
R3012 VSS.n421 VSS.n420 22.72
R3013 VSS.n419 VSS.n418 22.72
R3014 VSS.n417 VSS.n416 22.72
R3015 VSS.n415 VSS.n414 22.72
R3016 VSS.n343 VSS.n341 22.67
R3017 VSS.n344 VSS.n340 22.67
R3018 VSS.n345 VSS.n339 22.67
R3019 VSS.n346 VSS.n338 22.67
R3020 VSS.n347 VSS.n337 22.67
R3021 VSS.n348 VSS.n336 22.67
R3022 VSS.n349 VSS.n335 22.67
R3023 VSS.n333 VSS.n330 21.678
R3024 VSS.n1612 VSS.n1611 18.823
R3025 VSS.n1083 VSS.n1082 18.07
R3026 VSS.t978 VSS.t2360 12.446
R3027 VSS.t1481 VSS.t1010 12.446
R3028 VSS.t2034 VSS.t405 12.446
R3029 VSS.t2048 VSS.t1502 12.446
R3030 VSS.t921 VSS.t2068 12.446
R3031 VSS.t869 VSS.t863 12.446
R3032 VSS.t498 VSS.t1763 12.446
R3033 VSS.t1458 VSS.t1247 12.446
R3034 VSS.t1461 VSS.t972 12.446
R3035 VSS.t1565 VSS.t846 12.446
R3036 VSS.t2420 VSS.t2504 12.446
R3037 VSS.t1122 VSS.t1173 12.446
R3038 VSS.t399 VSS.t1783 12.446
R3039 VSS.t154 VSS.t801 12.446
R3040 VSS.t1930 VSS.t2512 12.446
R3041 VSS.t1464 VSS.t907 12.446
R3042 VSS.n2160 VSS.n2159 10.352
R3043 VSS.n1934 VSS.n1933 10.352
R3044 VSS.n571 VSS.n570 10.352
R3045 VSS.n2256 VSS.n2255 10.343
R3046 VSS.n2030 VSS.n2029 10.343
R3047 VSS.n780 VSS.n779 10.343
R3048 VSS.n684 VSS.n683 10.343
R3049 VSS.n475 VSS.n474 10.343
R3050 VSS.n459 VSS.n443 10.077
R3051 VSS.n2273 VSS.n2272 10.026
R3052 VSS.n4 VSS.n1 9.652
R3053 VSS.n194 VSS.n192 9.558
R3054 VSS.n137 VSS.t161 8.401
R3055 VSS.n128 VSS.t1023 8.401
R3056 VSS.n119 VSS.t2438 8.401
R3057 VSS.n110 VSS.t1926 8.401
R3058 VSS.n101 VSS.t1577 8.401
R3059 VSS.n92 VSS.t2458 8.401
R3060 VSS.n83 VSS.t1066 8.401
R3061 VSS.n74 VSS.t103 8.401
R3062 VSS.n65 VSS.t784 8.401
R3063 VSS.n56 VSS.t1211 8.401
R3064 VSS.n47 VSS.t1158 8.401
R3065 VSS.n38 VSS.t986 8.401
R3066 VSS.n29 VSS.t2134 8.401
R3067 VSS.n20 VSS.t2317 8.401
R3068 VSS.n11 VSS.t2100 8.401
R3069 VSS.n2 VSS.t1398 8.401
R3070 VSS.n5 VSS.t1400 8.401
R3071 VSS.n14 VSS.t2097 8.401
R3072 VSS.n23 VSS.t2314 8.401
R3073 VSS.n32 VSS.t2131 8.401
R3074 VSS.n41 VSS.t988 8.401
R3075 VSS.n50 VSS.t1155 8.401
R3076 VSS.n59 VSS.t1213 8.401
R3077 VSS.n68 VSS.t781 8.401
R3078 VSS.n77 VSS.t101 8.401
R3079 VSS.n86 VSS.t496 8.401
R3080 VSS.n95 VSS.t2455 8.401
R3081 VSS.n104 VSS.t1579 8.401
R3082 VSS.n113 VSS.t1928 8.401
R3083 VSS.n122 VSS.t2435 8.401
R3084 VSS.n131 VSS.t1025 8.401
R3085 VSS.n331 VSS.t92 8.401
R3086 VSS.n185 VSS.t3 8.401
R3087 VSS.n182 VSS.t1024 8.401
R3088 VSS.n179 VSS.t2439 8.401
R3089 VSS.n176 VSS.t1927 8.401
R3090 VSS.n173 VSS.t1578 8.401
R3091 VSS.n170 VSS.t2459 8.401
R3092 VSS.n167 VSS.t2194 8.401
R3093 VSS.n164 VSS.t100 8.401
R3094 VSS.n161 VSS.t785 8.401
R3095 VSS.n158 VSS.t1212 8.401
R3096 VSS.n155 VSS.t1159 8.401
R3097 VSS.n152 VSS.t987 8.401
R3098 VSS.n149 VSS.t2135 8.401
R3099 VSS.n146 VSS.t2318 8.401
R3100 VSS.n143 VSS.t2101 8.401
R3101 VSS.n140 VSS.t1399 8.401
R3102 VSS.n193 VSS.t1397 8.401
R3103 VSS.n202 VSS.t2099 8.401
R3104 VSS.n211 VSS.t2316 8.401
R3105 VSS.n220 VSS.t2133 8.401
R3106 VSS.n229 VSS.t985 8.401
R3107 VSS.n238 VSS.t1157 8.401
R3108 VSS.n247 VSS.t1210 8.401
R3109 VSS.n256 VSS.t783 8.401
R3110 VSS.n265 VSS.t102 8.401
R3111 VSS.n274 VSS.t1065 8.401
R3112 VSS.n283 VSS.t2457 8.401
R3113 VSS.n292 VSS.t1576 8.401
R3114 VSS.n301 VSS.t1925 8.401
R3115 VSS.n310 VSS.t2437 8.401
R3116 VSS.n319 VSS.t1022 8.401
R3117 VSS.n328 VSS.t93 8.401
R3118 VSS.n330 VSS.n186 8.292
R3119 VSS.n1084 VSS.n1083 8.28
R3120 VSS.n1613 VSS.n1612 8.28
R3121 VSS.n2097 VSS.n2096 8.28
R3122 VSS.n621 VSS.n620 8.28
R3123 VSS.n2335 VSS.n2334 7.996
R3124 VSS.n334 VSS.n333 6.955
R3125 VSS.n2338 VSS.n2337 6.48
R3126 VSS.n219 VSS.n212 6.433
R3127 VSS.n210 VSS.n203 6.433
R3128 VSS.n145 VSS.n144 6.419
R3129 VSS.n148 VSS.n147 6.419
R3130 VSS.n237 VSS.n230 6.406
R3131 VSS.n228 VSS.n221 6.406
R3132 VSS.n151 VSS.n150 6.392
R3133 VSS.n154 VSS.n153 6.392
R3134 VSS.n318 VSS.n311 6.388
R3135 VSS.n291 VSS.n284 6.388
R3136 VSS.n282 VSS.n275 6.388
R3137 VSS.n273 VSS.n266 6.388
R3138 VSS.n264 VSS.n257 6.388
R3139 VSS.n255 VSS.n248 6.388
R3140 VSS.n246 VSS.n239 6.388
R3141 VSS.n309 VSS.n302 6.38
R3142 VSS.n300 VSS.n293 6.38
R3143 VSS.n25 VSS.n24 6.38
R3144 VSS.n16 VSS.n15 6.38
R3145 VSS.n19 VSS.n13 6.38
R3146 VSS.n28 VSS.n22 6.38
R3147 VSS.n157 VSS.n156 6.374
R3148 VSS.n160 VSS.n159 6.374
R3149 VSS.n163 VSS.n162 6.374
R3150 VSS.n166 VSS.n165 6.374
R3151 VSS.n169 VSS.n168 6.374
R3152 VSS.n172 VSS.n171 6.374
R3153 VSS.n181 VSS.n180 6.374
R3154 VSS.n175 VSS.n174 6.366
R3155 VSS.n178 VSS.n177 6.366
R3156 VSS.n2335 VSS.n2288 6.36
R3157 VSS.n43 VSS.n42 6.354
R3158 VSS.n34 VSS.n33 6.354
R3159 VSS.n37 VSS.n31 6.353
R3160 VSS.n46 VSS.n40 6.353
R3161 VSS.n124 VSS.n123 6.336
R3162 VSS.n97 VSS.n96 6.336
R3163 VSS.n88 VSS.n87 6.336
R3164 VSS.n79 VSS.n78 6.336
R3165 VSS.n70 VSS.n69 6.336
R3166 VSS.n61 VSS.n60 6.336
R3167 VSS.n52 VSS.n51 6.336
R3168 VSS.n55 VSS.n49 6.335
R3169 VSS.n64 VSS.n58 6.335
R3170 VSS.n73 VSS.n67 6.335
R3171 VSS.n82 VSS.n76 6.335
R3172 VSS.n91 VSS.n85 6.335
R3173 VSS.n100 VSS.n94 6.335
R3174 VSS.n127 VSS.n121 6.335
R3175 VSS.n115 VSS.n114 6.327
R3176 VSS.n106 VSS.n105 6.327
R3177 VSS.n109 VSS.n103 6.326
R3178 VSS.n118 VSS.n112 6.326
R3179 VSS.n1710 VSS.n1709 6.299
R3180 VSS.n1565 VSS.n1564 6.299
R3181 VSS.n1181 VSS.n1180 6.299
R3182 VSS.n748 VSS.n747 6.299
R3183 VSS.n652 VSS.n651 6.299
R3184 VSS.n539 VSS.n538 6.299
R3185 VSS.n1998 VSS.n1997 6.291
R3186 VSS.n2288 VSS.n2287 6.29
R3187 VSS.n1838 VSS.n1837 6.29
R3188 VSS.n1501 VSS.n1500 6.29
R3189 VSS.n1437 VSS.n1436 6.29
R3190 VSS.n1373 VSS.n1372 6.29
R3191 VSS.n1309 VSS.n1308 6.29
R3192 VSS.n1245 VSS.n1244 6.29
R3193 VSS.n1036 VSS.n1035 6.29
R3194 VSS.n972 VSS.n971 6.29
R3195 VSS.n908 VSS.n907 6.29
R3196 VSS.n844 VSS.n843 6.29
R3197 VSS.n2128 VSS.n2127 6.29
R3198 VSS.n1646 VSS.n1645 6.29
R3199 VSS.n1117 VSS.n1116 6.29
R3200 VSS.n1774 VSS.n1773 6.281
R3201 VSS.n2224 VSS.n2223 6.276
R3202 VSS.n1902 VSS.n1901 6.276
R3203 VSS.t2355 VSS.t2084 6.223
R3204 VSS.t1280 VSS.t501 6.223
R3205 VSS.t395 VSS.t2033 6.223
R3206 VSS.t1352 VSS.t2177 6.223
R3207 VSS.t2115 VSS.t1827 6.223
R3208 VSS.t1699 VSS.t88 6.223
R3209 VSS.t2017 VSS.t1432 6.223
R3210 VSS.t1936 VSS.t1659 6.223
R3211 VSS.t1813 VSS.t45 6.223
R3212 VSS.t949 VSS.t1427 6.223
R3213 VSS.t445 VSS.t408 6.223
R3214 VSS.t1731 VSS.t1704 6.223
R3215 VSS.t1642 VSS.t1129 6.223
R3216 VSS.t1998 VSS.t2493 6.223
R3217 VSS.t1693 VSS.t1938 6.223
R3218 VSS.t1902 VSS.t937 6.223
R3219 VSS.n327 VSS.n320 6.103
R3220 VSS.n184 VSS.n183 6.089
R3221 VSS.n133 VSS.n132 6.05
R3222 VSS.n136 VSS.n130 6.049
R3223 VSS.n330 VSS.n329 5.835
R3224 VSS.n333 VSS.n332 5.835
R3225 VSS.n10 VSS.n9 5.702
R3226 VSS.n19 VSS.n18 5.702
R3227 VSS.n28 VSS.n27 5.702
R3228 VSS.n37 VSS.n36 5.702
R3229 VSS.n46 VSS.n45 5.702
R3230 VSS.n55 VSS.n54 5.702
R3231 VSS.n64 VSS.n63 5.702
R3232 VSS.n73 VSS.n72 5.702
R3233 VSS.n82 VSS.n81 5.702
R3234 VSS.n91 VSS.n90 5.702
R3235 VSS.n100 VSS.n99 5.702
R3236 VSS.n109 VSS.n108 5.702
R3237 VSS.n118 VSS.n117 5.702
R3238 VSS.n127 VSS.n126 5.702
R3239 VSS.n136 VSS.n135 5.702
R3240 VSS.n201 VSS.n200 5.662
R3241 VSS.n210 VSS.n209 5.662
R3242 VSS.n219 VSS.n218 5.662
R3243 VSS.n228 VSS.n227 5.662
R3244 VSS.n237 VSS.n236 5.662
R3245 VSS.n246 VSS.n245 5.662
R3246 VSS.n255 VSS.n254 5.662
R3247 VSS.n264 VSS.n263 5.662
R3248 VSS.n273 VSS.n272 5.662
R3249 VSS.n282 VSS.n281 5.662
R3250 VSS.n291 VSS.n290 5.662
R3251 VSS.n300 VSS.n299 5.662
R3252 VSS.n309 VSS.n308 5.662
R3253 VSS.n318 VSS.n317 5.662
R3254 VSS.n327 VSS.n326 5.662
R3255 VSS.n9 VSS.n7 5.615
R3256 VSS.n18 VSS.n16 5.615
R3257 VSS.n27 VSS.n25 5.615
R3258 VSS.n36 VSS.n34 5.615
R3259 VSS.n45 VSS.n43 5.615
R3260 VSS.n54 VSS.n52 5.615
R3261 VSS.n63 VSS.n61 5.615
R3262 VSS.n72 VSS.n70 5.615
R3263 VSS.n81 VSS.n79 5.615
R3264 VSS.n90 VSS.n88 5.615
R3265 VSS.n99 VSS.n97 5.615
R3266 VSS.n108 VSS.n106 5.615
R3267 VSS.n117 VSS.n115 5.615
R3268 VSS.n126 VSS.n124 5.615
R3269 VSS.n135 VSS.n133 5.615
R3270 VSS.n2336 VSS.n2335 5.536
R3271 VSS.n459 VSS.n458 5.416
R3272 VSS.n2144 VSS.n2143 5.409
R3273 VSS.n2240 VSS.n2239 5.407
R3274 VSS.n2014 VSS.n2013 5.407
R3275 VSS.n1918 VSS.n1917 5.407
R3276 VSS.n555 VSS.n554 5.407
R3277 VSS.n668 VSS.n667 5.4
R3278 VSS.n764 VSS.n763 5.398
R3279 VSS.n2274 VSS.n2273 5.133
R3280 VSS.n2275 VSS.n2274 5.133
R3281 VSS.n2276 VSS.n2275 5.133
R3282 VSS.n2277 VSS.n2276 5.133
R3283 VSS.n2278 VSS.n2277 5.133
R3284 VSS.n2279 VSS.n2278 5.133
R3285 VSS.n2280 VSS.n2279 5.133
R3286 VSS.n2281 VSS.n2280 5.133
R3287 VSS.n2282 VSS.n2281 5.133
R3288 VSS.n2283 VSS.n2282 5.133
R3289 VSS.n2284 VSS.n2283 5.133
R3290 VSS.n2285 VSS.n2284 5.133
R3291 VSS.n2286 VSS.n2285 5.133
R3292 VSS.n2287 VSS.n2286 5.133
R3293 VSS.n2130 VSS.n2129 4.999
R3294 VSS.n2131 VSS.n2130 4.999
R3295 VSS.n2132 VSS.n2131 4.999
R3296 VSS.n2133 VSS.n2132 4.999
R3297 VSS.n2134 VSS.n2133 4.999
R3298 VSS.n2135 VSS.n2134 4.999
R3299 VSS.n2136 VSS.n2135 4.999
R3300 VSS.n2137 VSS.n2136 4.999
R3301 VSS.n2138 VSS.n2137 4.999
R3302 VSS.n2139 VSS.n2138 4.999
R3303 VSS.n2140 VSS.n2139 4.999
R3304 VSS.n2141 VSS.n2140 4.999
R3305 VSS.n2142 VSS.n2141 4.999
R3306 VSS.n2143 VSS.n2142 4.999
R3307 VSS.n654 VSS.n653 4.999
R3308 VSS.n655 VSS.n654 4.999
R3309 VSS.n656 VSS.n655 4.999
R3310 VSS.n657 VSS.n656 4.999
R3311 VSS.n658 VSS.n657 4.999
R3312 VSS.n659 VSS.n658 4.999
R3313 VSS.n660 VSS.n659 4.999
R3314 VSS.n661 VSS.n660 4.999
R3315 VSS.n662 VSS.n661 4.999
R3316 VSS.n663 VSS.n662 4.999
R3317 VSS.n664 VSS.n663 4.999
R3318 VSS.n665 VSS.n664 4.999
R3319 VSS.n666 VSS.n665 4.999
R3320 VSS.n667 VSS.n666 4.999
R3321 VSS.n2226 VSS.n2225 4.994
R3322 VSS.n2227 VSS.n2226 4.994
R3323 VSS.n2228 VSS.n2227 4.994
R3324 VSS.n2229 VSS.n2228 4.994
R3325 VSS.n2230 VSS.n2229 4.994
R3326 VSS.n2231 VSS.n2230 4.994
R3327 VSS.n2232 VSS.n2231 4.994
R3328 VSS.n2233 VSS.n2232 4.994
R3329 VSS.n2234 VSS.n2233 4.994
R3330 VSS.n2235 VSS.n2234 4.994
R3331 VSS.n2236 VSS.n2235 4.994
R3332 VSS.n2237 VSS.n2236 4.994
R3333 VSS.n2238 VSS.n2237 4.994
R3334 VSS.n2239 VSS.n2238 4.994
R3335 VSS.n2000 VSS.n1999 4.994
R3336 VSS.n2001 VSS.n2000 4.994
R3337 VSS.n2002 VSS.n2001 4.994
R3338 VSS.n2003 VSS.n2002 4.994
R3339 VSS.n2004 VSS.n2003 4.994
R3340 VSS.n2005 VSS.n2004 4.994
R3341 VSS.n2006 VSS.n2005 4.994
R3342 VSS.n2007 VSS.n2006 4.994
R3343 VSS.n2008 VSS.n2007 4.994
R3344 VSS.n2009 VSS.n2008 4.994
R3345 VSS.n2010 VSS.n2009 4.994
R3346 VSS.n2011 VSS.n2010 4.994
R3347 VSS.n2012 VSS.n2011 4.994
R3348 VSS.n2013 VSS.n2012 4.994
R3349 VSS.n1904 VSS.n1903 4.994
R3350 VSS.n1905 VSS.n1904 4.994
R3351 VSS.n1906 VSS.n1905 4.994
R3352 VSS.n1907 VSS.n1906 4.994
R3353 VSS.n1908 VSS.n1907 4.994
R3354 VSS.n1909 VSS.n1908 4.994
R3355 VSS.n1910 VSS.n1909 4.994
R3356 VSS.n1911 VSS.n1910 4.994
R3357 VSS.n1912 VSS.n1911 4.994
R3358 VSS.n1913 VSS.n1912 4.994
R3359 VSS.n1914 VSS.n1913 4.994
R3360 VSS.n1915 VSS.n1914 4.994
R3361 VSS.n1916 VSS.n1915 4.994
R3362 VSS.n1917 VSS.n1916 4.994
R3363 VSS.n750 VSS.n749 4.994
R3364 VSS.n751 VSS.n750 4.994
R3365 VSS.n752 VSS.n751 4.994
R3366 VSS.n753 VSS.n752 4.994
R3367 VSS.n754 VSS.n753 4.994
R3368 VSS.n755 VSS.n754 4.994
R3369 VSS.n756 VSS.n755 4.994
R3370 VSS.n757 VSS.n756 4.994
R3371 VSS.n758 VSS.n757 4.994
R3372 VSS.n759 VSS.n758 4.994
R3373 VSS.n760 VSS.n759 4.994
R3374 VSS.n761 VSS.n760 4.994
R3375 VSS.n762 VSS.n761 4.994
R3376 VSS.n763 VSS.n762 4.994
R3377 VSS.n541 VSS.n540 4.994
R3378 VSS.n542 VSS.n541 4.994
R3379 VSS.n543 VSS.n542 4.994
R3380 VSS.n544 VSS.n543 4.994
R3381 VSS.n545 VSS.n544 4.994
R3382 VSS.n546 VSS.n545 4.994
R3383 VSS.n547 VSS.n546 4.994
R3384 VSS.n548 VSS.n547 4.994
R3385 VSS.n549 VSS.n548 4.994
R3386 VSS.n550 VSS.n549 4.994
R3387 VSS.n551 VSS.n550 4.994
R3388 VSS.n552 VSS.n551 4.994
R3389 VSS.n553 VSS.n552 4.994
R3390 VSS.n554 VSS.n553 4.994
R3391 VSS.n445 VSS.n444 4.994
R3392 VSS.n446 VSS.n445 4.994
R3393 VSS.n447 VSS.n446 4.994
R3394 VSS.n448 VSS.n447 4.994
R3395 VSS.n449 VSS.n448 4.994
R3396 VSS.n450 VSS.n449 4.994
R3397 VSS.n451 VSS.n450 4.994
R3398 VSS.n452 VSS.n451 4.994
R3399 VSS.n453 VSS.n452 4.994
R3400 VSS.n454 VSS.n453 4.994
R3401 VSS.n455 VSS.n454 4.994
R3402 VSS.n456 VSS.n455 4.994
R3403 VSS.n457 VSS.n456 4.994
R3404 VSS.n458 VSS.n457 4.994
R3405 VSS.n2242 VSS.n2241 4.979
R3406 VSS.n2243 VSS.n2242 4.979
R3407 VSS.n2244 VSS.n2243 4.979
R3408 VSS.n2245 VSS.n2244 4.979
R3409 VSS.n2246 VSS.n2245 4.979
R3410 VSS.n2247 VSS.n2246 4.979
R3411 VSS.n2248 VSS.n2247 4.979
R3412 VSS.n2249 VSS.n2248 4.979
R3413 VSS.n2250 VSS.n2249 4.979
R3414 VSS.n2251 VSS.n2250 4.979
R3415 VSS.n2252 VSS.n2251 4.979
R3416 VSS.n2253 VSS.n2252 4.979
R3417 VSS.n2254 VSS.n2253 4.979
R3418 VSS.n2255 VSS.n2254 4.979
R3419 VSS.n2146 VSS.n2145 4.979
R3420 VSS.n2147 VSS.n2146 4.979
R3421 VSS.n2148 VSS.n2147 4.979
R3422 VSS.n2149 VSS.n2148 4.979
R3423 VSS.n2150 VSS.n2149 4.979
R3424 VSS.n2151 VSS.n2150 4.979
R3425 VSS.n2152 VSS.n2151 4.979
R3426 VSS.n2153 VSS.n2152 4.979
R3427 VSS.n2154 VSS.n2153 4.979
R3428 VSS.n2155 VSS.n2154 4.979
R3429 VSS.n2156 VSS.n2155 4.979
R3430 VSS.n2157 VSS.n2156 4.979
R3431 VSS.n2158 VSS.n2157 4.979
R3432 VSS.n2159 VSS.n2158 4.979
R3433 VSS.n2016 VSS.n2015 4.979
R3434 VSS.n2017 VSS.n2016 4.979
R3435 VSS.n2018 VSS.n2017 4.979
R3436 VSS.n2019 VSS.n2018 4.979
R3437 VSS.n2020 VSS.n2019 4.979
R3438 VSS.n2021 VSS.n2020 4.979
R3439 VSS.n2022 VSS.n2021 4.979
R3440 VSS.n2023 VSS.n2022 4.979
R3441 VSS.n2024 VSS.n2023 4.979
R3442 VSS.n2025 VSS.n2024 4.979
R3443 VSS.n2026 VSS.n2025 4.979
R3444 VSS.n2027 VSS.n2026 4.979
R3445 VSS.n2028 VSS.n2027 4.979
R3446 VSS.n2029 VSS.n2028 4.979
R3447 VSS.n1920 VSS.n1919 4.979
R3448 VSS.n1921 VSS.n1920 4.979
R3449 VSS.n1922 VSS.n1921 4.979
R3450 VSS.n1923 VSS.n1922 4.979
R3451 VSS.n1924 VSS.n1923 4.979
R3452 VSS.n1925 VSS.n1924 4.979
R3453 VSS.n1926 VSS.n1925 4.979
R3454 VSS.n1927 VSS.n1926 4.979
R3455 VSS.n1928 VSS.n1927 4.979
R3456 VSS.n1929 VSS.n1928 4.979
R3457 VSS.n1930 VSS.n1929 4.979
R3458 VSS.n1931 VSS.n1930 4.979
R3459 VSS.n1932 VSS.n1931 4.979
R3460 VSS.n1933 VSS.n1932 4.979
R3461 VSS.n766 VSS.n765 4.979
R3462 VSS.n767 VSS.n766 4.979
R3463 VSS.n768 VSS.n767 4.979
R3464 VSS.n769 VSS.n768 4.979
R3465 VSS.n770 VSS.n769 4.979
R3466 VSS.n771 VSS.n770 4.979
R3467 VSS.n772 VSS.n771 4.979
R3468 VSS.n773 VSS.n772 4.979
R3469 VSS.n774 VSS.n773 4.979
R3470 VSS.n775 VSS.n774 4.979
R3471 VSS.n776 VSS.n775 4.979
R3472 VSS.n777 VSS.n776 4.979
R3473 VSS.n778 VSS.n777 4.979
R3474 VSS.n779 VSS.n778 4.979
R3475 VSS.n670 VSS.n669 4.979
R3476 VSS.n671 VSS.n670 4.979
R3477 VSS.n672 VSS.n671 4.979
R3478 VSS.n673 VSS.n672 4.979
R3479 VSS.n674 VSS.n673 4.979
R3480 VSS.n675 VSS.n674 4.979
R3481 VSS.n676 VSS.n675 4.979
R3482 VSS.n677 VSS.n676 4.979
R3483 VSS.n678 VSS.n677 4.979
R3484 VSS.n679 VSS.n678 4.979
R3485 VSS.n680 VSS.n679 4.979
R3486 VSS.n681 VSS.n680 4.979
R3487 VSS.n682 VSS.n681 4.979
R3488 VSS.n683 VSS.n682 4.979
R3489 VSS.n557 VSS.n556 4.979
R3490 VSS.n558 VSS.n557 4.979
R3491 VSS.n559 VSS.n558 4.979
R3492 VSS.n560 VSS.n559 4.979
R3493 VSS.n561 VSS.n560 4.979
R3494 VSS.n562 VSS.n561 4.979
R3495 VSS.n563 VSS.n562 4.979
R3496 VSS.n564 VSS.n563 4.979
R3497 VSS.n565 VSS.n564 4.979
R3498 VSS.n566 VSS.n565 4.979
R3499 VSS.n567 VSS.n566 4.979
R3500 VSS.n568 VSS.n567 4.979
R3501 VSS.n569 VSS.n568 4.979
R3502 VSS.n570 VSS.n569 4.979
R3503 VSS.n461 VSS.n460 4.979
R3504 VSS.n462 VSS.n461 4.979
R3505 VSS.n463 VSS.n462 4.979
R3506 VSS.n464 VSS.n463 4.979
R3507 VSS.n465 VSS.n464 4.979
R3508 VSS.n466 VSS.n465 4.979
R3509 VSS.n467 VSS.n466 4.979
R3510 VSS.n468 VSS.n467 4.979
R3511 VSS.n469 VSS.n468 4.979
R3512 VSS.n470 VSS.n469 4.979
R3513 VSS.n471 VSS.n470 4.979
R3514 VSS.n472 VSS.n471 4.979
R3515 VSS.n473 VSS.n472 4.979
R3516 VSS.n474 VSS.n473 4.979
R3517 VSS.n417 VSS.n415 4.97
R3518 VSS.n419 VSS.n417 4.97
R3519 VSS.n421 VSS.n419 4.97
R3520 VSS.n423 VSS.n421 4.97
R3521 VSS.n425 VSS.n423 4.97
R3522 VSS.n427 VSS.n425 4.97
R3523 VSS.n429 VSS.n427 4.97
R3524 VSS.n431 VSS.n429 4.97
R3525 VSS.n433 VSS.n431 4.97
R3526 VSS.n435 VSS.n433 4.97
R3527 VSS.n437 VSS.n435 4.97
R3528 VSS.n439 VSS.n437 4.97
R3529 VSS.n441 VSS.n439 4.97
R3530 VSS.n443 VSS.n441 4.97
R3531 VSS.n2273 VSS.n2271 4.893
R3532 VSS.n2274 VSS.n2270 4.893
R3533 VSS.n2275 VSS.n2269 4.893
R3534 VSS.n2276 VSS.n2268 4.893
R3535 VSS.n2277 VSS.n2267 4.893
R3536 VSS.n2278 VSS.n2266 4.893
R3537 VSS.n2279 VSS.n2265 4.893
R3538 VSS.n2280 VSS.n2264 4.893
R3539 VSS.n2281 VSS.n2263 4.893
R3540 VSS.n2282 VSS.n2262 4.893
R3541 VSS.n2283 VSS.n2261 4.893
R3542 VSS.n2284 VSS.n2260 4.893
R3543 VSS.n2285 VSS.n2259 4.893
R3544 VSS.n2286 VSS.n2258 4.893
R3545 VSS.n2287 VSS.n2257 4.893
R3546 VSS.n2178 VSS.n2176 4.893
R3547 VSS.n2181 VSS.n2175 4.893
R3548 VSS.n2184 VSS.n2174 4.893
R3549 VSS.n2187 VSS.n2173 4.893
R3550 VSS.n2190 VSS.n2172 4.893
R3551 VSS.n2193 VSS.n2171 4.893
R3552 VSS.n2196 VSS.n2170 4.893
R3553 VSS.n2199 VSS.n2169 4.893
R3554 VSS.n2202 VSS.n2168 4.893
R3555 VSS.n2205 VSS.n2167 4.893
R3556 VSS.n2208 VSS.n2166 4.893
R3557 VSS.n2211 VSS.n2165 4.893
R3558 VSS.n2214 VSS.n2164 4.893
R3559 VSS.n2217 VSS.n2163 4.893
R3560 VSS.n2220 VSS.n2162 4.893
R3561 VSS.n2223 VSS.n2161 4.893
R3562 VSS.n1952 VSS.n1950 4.893
R3563 VSS.n1955 VSS.n1949 4.893
R3564 VSS.n1958 VSS.n1948 4.893
R3565 VSS.n1961 VSS.n1947 4.893
R3566 VSS.n1964 VSS.n1946 4.893
R3567 VSS.n1967 VSS.n1945 4.893
R3568 VSS.n1970 VSS.n1944 4.893
R3569 VSS.n1973 VSS.n1943 4.893
R3570 VSS.n1976 VSS.n1942 4.893
R3571 VSS.n1979 VSS.n1941 4.893
R3572 VSS.n1982 VSS.n1940 4.893
R3573 VSS.n1985 VSS.n1939 4.893
R3574 VSS.n1988 VSS.n1938 4.893
R3575 VSS.n1991 VSS.n1937 4.893
R3576 VSS.n1994 VSS.n1936 4.893
R3577 VSS.n1997 VSS.n1935 4.893
R3578 VSS.n1856 VSS.n1854 4.893
R3579 VSS.n1859 VSS.n1853 4.893
R3580 VSS.n1862 VSS.n1852 4.893
R3581 VSS.n1865 VSS.n1851 4.893
R3582 VSS.n1868 VSS.n1850 4.893
R3583 VSS.n1871 VSS.n1849 4.893
R3584 VSS.n1874 VSS.n1848 4.893
R3585 VSS.n1877 VSS.n1847 4.893
R3586 VSS.n1880 VSS.n1846 4.893
R3587 VSS.n1883 VSS.n1845 4.893
R3588 VSS.n1886 VSS.n1844 4.893
R3589 VSS.n1889 VSS.n1843 4.893
R3590 VSS.n1892 VSS.n1842 4.893
R3591 VSS.n1895 VSS.n1841 4.893
R3592 VSS.n1898 VSS.n1840 4.893
R3593 VSS.n1901 VSS.n1839 4.893
R3594 VSS.n1792 VSS.n1790 4.893
R3595 VSS.n1795 VSS.n1789 4.893
R3596 VSS.n1798 VSS.n1788 4.893
R3597 VSS.n1801 VSS.n1787 4.893
R3598 VSS.n1804 VSS.n1786 4.893
R3599 VSS.n1807 VSS.n1785 4.893
R3600 VSS.n1810 VSS.n1784 4.893
R3601 VSS.n1813 VSS.n1783 4.893
R3602 VSS.n1816 VSS.n1782 4.893
R3603 VSS.n1819 VSS.n1781 4.893
R3604 VSS.n1822 VSS.n1780 4.893
R3605 VSS.n1825 VSS.n1779 4.893
R3606 VSS.n1828 VSS.n1778 4.893
R3607 VSS.n1831 VSS.n1777 4.893
R3608 VSS.n1834 VSS.n1776 4.893
R3609 VSS.n1837 VSS.n1775 4.893
R3610 VSS.n1728 VSS.n1726 4.893
R3611 VSS.n1731 VSS.n1725 4.893
R3612 VSS.n1734 VSS.n1724 4.893
R3613 VSS.n1737 VSS.n1723 4.893
R3614 VSS.n1740 VSS.n1722 4.893
R3615 VSS.n1743 VSS.n1721 4.893
R3616 VSS.n1746 VSS.n1720 4.893
R3617 VSS.n1749 VSS.n1719 4.893
R3618 VSS.n1752 VSS.n1718 4.893
R3619 VSS.n1755 VSS.n1717 4.893
R3620 VSS.n1758 VSS.n1716 4.893
R3621 VSS.n1761 VSS.n1715 4.893
R3622 VSS.n1764 VSS.n1714 4.893
R3623 VSS.n1767 VSS.n1713 4.893
R3624 VSS.n1770 VSS.n1712 4.893
R3625 VSS.n1773 VSS.n1711 4.893
R3626 VSS.n1664 VSS.n1662 4.893
R3627 VSS.n1667 VSS.n1661 4.893
R3628 VSS.n1670 VSS.n1660 4.893
R3629 VSS.n1673 VSS.n1659 4.893
R3630 VSS.n1676 VSS.n1658 4.893
R3631 VSS.n1679 VSS.n1657 4.893
R3632 VSS.n1682 VSS.n1656 4.893
R3633 VSS.n1685 VSS.n1655 4.893
R3634 VSS.n1688 VSS.n1654 4.893
R3635 VSS.n1691 VSS.n1653 4.893
R3636 VSS.n1694 VSS.n1652 4.893
R3637 VSS.n1697 VSS.n1651 4.893
R3638 VSS.n1700 VSS.n1650 4.893
R3639 VSS.n1703 VSS.n1649 4.893
R3640 VSS.n1706 VSS.n1648 4.893
R3641 VSS.n1709 VSS.n1647 4.893
R3642 VSS.n1519 VSS.n1517 4.893
R3643 VSS.n1522 VSS.n1516 4.893
R3644 VSS.n1525 VSS.n1515 4.893
R3645 VSS.n1528 VSS.n1514 4.893
R3646 VSS.n1531 VSS.n1513 4.893
R3647 VSS.n1534 VSS.n1512 4.893
R3648 VSS.n1537 VSS.n1511 4.893
R3649 VSS.n1540 VSS.n1510 4.893
R3650 VSS.n1543 VSS.n1509 4.893
R3651 VSS.n1546 VSS.n1508 4.893
R3652 VSS.n1549 VSS.n1507 4.893
R3653 VSS.n1552 VSS.n1506 4.893
R3654 VSS.n1555 VSS.n1505 4.893
R3655 VSS.n1558 VSS.n1504 4.893
R3656 VSS.n1561 VSS.n1503 4.893
R3657 VSS.n1564 VSS.n1502 4.893
R3658 VSS.n1455 VSS.n1453 4.893
R3659 VSS.n1458 VSS.n1452 4.893
R3660 VSS.n1461 VSS.n1451 4.893
R3661 VSS.n1464 VSS.n1450 4.893
R3662 VSS.n1467 VSS.n1449 4.893
R3663 VSS.n1470 VSS.n1448 4.893
R3664 VSS.n1473 VSS.n1447 4.893
R3665 VSS.n1476 VSS.n1446 4.893
R3666 VSS.n1479 VSS.n1445 4.893
R3667 VSS.n1482 VSS.n1444 4.893
R3668 VSS.n1485 VSS.n1443 4.893
R3669 VSS.n1488 VSS.n1442 4.893
R3670 VSS.n1491 VSS.n1441 4.893
R3671 VSS.n1494 VSS.n1440 4.893
R3672 VSS.n1497 VSS.n1439 4.893
R3673 VSS.n1500 VSS.n1438 4.893
R3674 VSS.n1391 VSS.n1389 4.893
R3675 VSS.n1394 VSS.n1388 4.893
R3676 VSS.n1397 VSS.n1387 4.893
R3677 VSS.n1400 VSS.n1386 4.893
R3678 VSS.n1403 VSS.n1385 4.893
R3679 VSS.n1406 VSS.n1384 4.893
R3680 VSS.n1409 VSS.n1383 4.893
R3681 VSS.n1412 VSS.n1382 4.893
R3682 VSS.n1415 VSS.n1381 4.893
R3683 VSS.n1418 VSS.n1380 4.893
R3684 VSS.n1421 VSS.n1379 4.893
R3685 VSS.n1424 VSS.n1378 4.893
R3686 VSS.n1427 VSS.n1377 4.893
R3687 VSS.n1430 VSS.n1376 4.893
R3688 VSS.n1433 VSS.n1375 4.893
R3689 VSS.n1436 VSS.n1374 4.893
R3690 VSS.n1327 VSS.n1325 4.893
R3691 VSS.n1330 VSS.n1324 4.893
R3692 VSS.n1333 VSS.n1323 4.893
R3693 VSS.n1336 VSS.n1322 4.893
R3694 VSS.n1339 VSS.n1321 4.893
R3695 VSS.n1342 VSS.n1320 4.893
R3696 VSS.n1345 VSS.n1319 4.893
R3697 VSS.n1348 VSS.n1318 4.893
R3698 VSS.n1351 VSS.n1317 4.893
R3699 VSS.n1354 VSS.n1316 4.893
R3700 VSS.n1357 VSS.n1315 4.893
R3701 VSS.n1360 VSS.n1314 4.893
R3702 VSS.n1363 VSS.n1313 4.893
R3703 VSS.n1366 VSS.n1312 4.893
R3704 VSS.n1369 VSS.n1311 4.893
R3705 VSS.n1372 VSS.n1310 4.893
R3706 VSS.n1263 VSS.n1261 4.893
R3707 VSS.n1266 VSS.n1260 4.893
R3708 VSS.n1269 VSS.n1259 4.893
R3709 VSS.n1272 VSS.n1258 4.893
R3710 VSS.n1275 VSS.n1257 4.893
R3711 VSS.n1278 VSS.n1256 4.893
R3712 VSS.n1281 VSS.n1255 4.893
R3713 VSS.n1284 VSS.n1254 4.893
R3714 VSS.n1287 VSS.n1253 4.893
R3715 VSS.n1290 VSS.n1252 4.893
R3716 VSS.n1293 VSS.n1251 4.893
R3717 VSS.n1296 VSS.n1250 4.893
R3718 VSS.n1299 VSS.n1249 4.893
R3719 VSS.n1302 VSS.n1248 4.893
R3720 VSS.n1305 VSS.n1247 4.893
R3721 VSS.n1308 VSS.n1246 4.893
R3722 VSS.n1199 VSS.n1197 4.893
R3723 VSS.n1202 VSS.n1196 4.893
R3724 VSS.n1205 VSS.n1195 4.893
R3725 VSS.n1208 VSS.n1194 4.893
R3726 VSS.n1211 VSS.n1193 4.893
R3727 VSS.n1214 VSS.n1192 4.893
R3728 VSS.n1217 VSS.n1191 4.893
R3729 VSS.n1220 VSS.n1190 4.893
R3730 VSS.n1223 VSS.n1189 4.893
R3731 VSS.n1226 VSS.n1188 4.893
R3732 VSS.n1229 VSS.n1187 4.893
R3733 VSS.n1232 VSS.n1186 4.893
R3734 VSS.n1235 VSS.n1185 4.893
R3735 VSS.n1238 VSS.n1184 4.893
R3736 VSS.n1241 VSS.n1183 4.893
R3737 VSS.n1244 VSS.n1182 4.893
R3738 VSS.n1135 VSS.n1133 4.893
R3739 VSS.n1138 VSS.n1132 4.893
R3740 VSS.n1141 VSS.n1131 4.893
R3741 VSS.n1144 VSS.n1130 4.893
R3742 VSS.n1147 VSS.n1129 4.893
R3743 VSS.n1150 VSS.n1128 4.893
R3744 VSS.n1153 VSS.n1127 4.893
R3745 VSS.n1156 VSS.n1126 4.893
R3746 VSS.n1159 VSS.n1125 4.893
R3747 VSS.n1162 VSS.n1124 4.893
R3748 VSS.n1165 VSS.n1123 4.893
R3749 VSS.n1168 VSS.n1122 4.893
R3750 VSS.n1171 VSS.n1121 4.893
R3751 VSS.n1174 VSS.n1120 4.893
R3752 VSS.n1177 VSS.n1119 4.893
R3753 VSS.n1180 VSS.n1118 4.893
R3754 VSS.n990 VSS.n988 4.893
R3755 VSS.n993 VSS.n987 4.893
R3756 VSS.n996 VSS.n986 4.893
R3757 VSS.n999 VSS.n985 4.893
R3758 VSS.n1002 VSS.n984 4.893
R3759 VSS.n1005 VSS.n983 4.893
R3760 VSS.n1008 VSS.n982 4.893
R3761 VSS.n1011 VSS.n981 4.893
R3762 VSS.n1014 VSS.n980 4.893
R3763 VSS.n1017 VSS.n979 4.893
R3764 VSS.n1020 VSS.n978 4.893
R3765 VSS.n1023 VSS.n977 4.893
R3766 VSS.n1026 VSS.n976 4.893
R3767 VSS.n1029 VSS.n975 4.893
R3768 VSS.n1032 VSS.n974 4.893
R3769 VSS.n1035 VSS.n973 4.893
R3770 VSS.n926 VSS.n924 4.893
R3771 VSS.n929 VSS.n923 4.893
R3772 VSS.n932 VSS.n922 4.893
R3773 VSS.n935 VSS.n921 4.893
R3774 VSS.n938 VSS.n920 4.893
R3775 VSS.n941 VSS.n919 4.893
R3776 VSS.n944 VSS.n918 4.893
R3777 VSS.n947 VSS.n917 4.893
R3778 VSS.n950 VSS.n916 4.893
R3779 VSS.n953 VSS.n915 4.893
R3780 VSS.n956 VSS.n914 4.893
R3781 VSS.n959 VSS.n913 4.893
R3782 VSS.n962 VSS.n912 4.893
R3783 VSS.n965 VSS.n911 4.893
R3784 VSS.n968 VSS.n910 4.893
R3785 VSS.n971 VSS.n909 4.893
R3786 VSS.n862 VSS.n860 4.893
R3787 VSS.n865 VSS.n859 4.893
R3788 VSS.n868 VSS.n858 4.893
R3789 VSS.n871 VSS.n857 4.893
R3790 VSS.n874 VSS.n856 4.893
R3791 VSS.n877 VSS.n855 4.893
R3792 VSS.n880 VSS.n854 4.893
R3793 VSS.n883 VSS.n853 4.893
R3794 VSS.n886 VSS.n852 4.893
R3795 VSS.n889 VSS.n851 4.893
R3796 VSS.n892 VSS.n850 4.893
R3797 VSS.n895 VSS.n849 4.893
R3798 VSS.n898 VSS.n848 4.893
R3799 VSS.n901 VSS.n847 4.893
R3800 VSS.n904 VSS.n846 4.893
R3801 VSS.n907 VSS.n845 4.893
R3802 VSS.n798 VSS.n796 4.893
R3803 VSS.n801 VSS.n795 4.893
R3804 VSS.n804 VSS.n794 4.893
R3805 VSS.n807 VSS.n793 4.893
R3806 VSS.n810 VSS.n792 4.893
R3807 VSS.n813 VSS.n791 4.893
R3808 VSS.n816 VSS.n790 4.893
R3809 VSS.n819 VSS.n789 4.893
R3810 VSS.n822 VSS.n788 4.893
R3811 VSS.n825 VSS.n787 4.893
R3812 VSS.n828 VSS.n786 4.893
R3813 VSS.n831 VSS.n785 4.893
R3814 VSS.n834 VSS.n784 4.893
R3815 VSS.n837 VSS.n783 4.893
R3816 VSS.n840 VSS.n782 4.893
R3817 VSS.n843 VSS.n781 4.893
R3818 VSS.n702 VSS.n700 4.893
R3819 VSS.n705 VSS.n699 4.893
R3820 VSS.n708 VSS.n698 4.893
R3821 VSS.n711 VSS.n697 4.893
R3822 VSS.n714 VSS.n696 4.893
R3823 VSS.n717 VSS.n695 4.893
R3824 VSS.n720 VSS.n694 4.893
R3825 VSS.n723 VSS.n693 4.893
R3826 VSS.n726 VSS.n692 4.893
R3827 VSS.n729 VSS.n691 4.893
R3828 VSS.n732 VSS.n690 4.893
R3829 VSS.n735 VSS.n689 4.893
R3830 VSS.n738 VSS.n688 4.893
R3831 VSS.n741 VSS.n687 4.893
R3832 VSS.n744 VSS.n686 4.893
R3833 VSS.n747 VSS.n685 4.893
R3834 VSS.n651 VSS.n573 4.893
R3835 VSS.n649 VSS.n576 4.893
R3836 VSS.n621 VSS.n618 4.893
R3837 VSS.n1613 VSS.n1610 4.893
R3838 VSS.n2097 VSS.n2093 4.893
R3839 VSS.n1084 VSS.n1081 4.893
R3840 VSS.n623 VSS.n615 4.893
R3841 VSS.n1615 VSS.n1607 4.893
R3842 VSS.n2099 VSS.n2089 4.893
R3843 VSS.n1086 VSS.n1078 4.893
R3844 VSS.n625 VSS.n612 4.893
R3845 VSS.n1617 VSS.n1604 4.893
R3846 VSS.n2101 VSS.n2085 4.893
R3847 VSS.n1088 VSS.n1075 4.893
R3848 VSS.n627 VSS.n609 4.893
R3849 VSS.n1619 VSS.n1601 4.893
R3850 VSS.n2103 VSS.n2081 4.893
R3851 VSS.n1090 VSS.n1072 4.893
R3852 VSS.n629 VSS.n606 4.893
R3853 VSS.n1621 VSS.n1598 4.893
R3854 VSS.n2105 VSS.n2077 4.893
R3855 VSS.n1092 VSS.n1069 4.893
R3856 VSS.n631 VSS.n603 4.893
R3857 VSS.n1623 VSS.n1595 4.893
R3858 VSS.n2107 VSS.n2073 4.893
R3859 VSS.n1094 VSS.n1066 4.893
R3860 VSS.n633 VSS.n600 4.893
R3861 VSS.n1625 VSS.n1592 4.893
R3862 VSS.n2109 VSS.n2069 4.893
R3863 VSS.n1096 VSS.n1063 4.893
R3864 VSS.n635 VSS.n597 4.893
R3865 VSS.n1627 VSS.n1589 4.893
R3866 VSS.n2111 VSS.n2065 4.893
R3867 VSS.n1098 VSS.n1060 4.893
R3868 VSS.n637 VSS.n594 4.893
R3869 VSS.n1629 VSS.n1586 4.893
R3870 VSS.n2113 VSS.n2061 4.893
R3871 VSS.n1100 VSS.n1057 4.893
R3872 VSS.n639 VSS.n591 4.893
R3873 VSS.n1631 VSS.n1583 4.893
R3874 VSS.n2115 VSS.n2057 4.893
R3875 VSS.n1102 VSS.n1054 4.893
R3876 VSS.n641 VSS.n588 4.893
R3877 VSS.n1633 VSS.n1580 4.893
R3878 VSS.n2117 VSS.n2053 4.893
R3879 VSS.n1104 VSS.n1051 4.893
R3880 VSS.n643 VSS.n585 4.893
R3881 VSS.n1635 VSS.n1577 4.893
R3882 VSS.n2119 VSS.n2049 4.893
R3883 VSS.n1106 VSS.n1048 4.893
R3884 VSS.n645 VSS.n582 4.893
R3885 VSS.n1637 VSS.n1574 4.893
R3886 VSS.n2121 VSS.n2045 4.893
R3887 VSS.n1108 VSS.n1045 4.893
R3888 VSS.n647 VSS.n579 4.893
R3889 VSS.n1639 VSS.n1571 4.893
R3890 VSS.n2123 VSS.n2041 4.893
R3891 VSS.n1110 VSS.n1042 4.893
R3892 VSS.n1116 VSS.n1038 4.893
R3893 VSS.n1114 VSS.n1113 4.893
R3894 VSS.n2125 VSS.n2037 4.893
R3895 VSS.n1641 VSS.n1568 4.893
R3896 VSS.n1645 VSS.n1644 4.893
R3897 VSS.n2127 VSS.n2033 4.893
R3898 VSS.n493 VSS.n491 4.893
R3899 VSS.n496 VSS.n490 4.893
R3900 VSS.n499 VSS.n489 4.893
R3901 VSS.n502 VSS.n488 4.893
R3902 VSS.n505 VSS.n487 4.893
R3903 VSS.n508 VSS.n486 4.893
R3904 VSS.n511 VSS.n485 4.893
R3905 VSS.n514 VSS.n484 4.893
R3906 VSS.n517 VSS.n483 4.893
R3907 VSS.n520 VSS.n482 4.893
R3908 VSS.n523 VSS.n481 4.893
R3909 VSS.n526 VSS.n480 4.893
R3910 VSS.n529 VSS.n479 4.893
R3911 VSS.n532 VSS.n478 4.893
R3912 VSS.n535 VSS.n477 4.893
R3913 VSS.n538 VSS.n476 4.893
R3914 VSS.n13 VSS.n10 3.95
R3915 VSS.n22 VSS.n19 3.95
R3916 VSS.n31 VSS.n28 3.95
R3917 VSS.n40 VSS.n37 3.95
R3918 VSS.n49 VSS.n46 3.95
R3919 VSS.n58 VSS.n55 3.95
R3920 VSS.n67 VSS.n64 3.95
R3921 VSS.n76 VSS.n73 3.95
R3922 VSS.n85 VSS.n82 3.95
R3923 VSS.n94 VSS.n91 3.95
R3924 VSS.n103 VSS.n100 3.95
R3925 VSS.n112 VSS.n109 3.95
R3926 VSS.n121 VSS.n118 3.95
R3927 VSS.n130 VSS.n127 3.95
R3928 VSS.n139 VSS.n136 3.95
R3929 VSS.n329 VSS.n327 3.896
R3930 VSS.n320 VSS.n318 3.896
R3931 VSS.n311 VSS.n309 3.896
R3932 VSS.n302 VSS.n300 3.896
R3933 VSS.n293 VSS.n291 3.896
R3934 VSS.n284 VSS.n282 3.896
R3935 VSS.n275 VSS.n273 3.896
R3936 VSS.n266 VSS.n264 3.896
R3937 VSS.n257 VSS.n255 3.896
R3938 VSS.n248 VSS.n246 3.896
R3939 VSS.n239 VSS.n237 3.896
R3940 VSS.n230 VSS.n228 3.896
R3941 VSS.n221 VSS.n219 3.896
R3942 VSS.n212 VSS.n210 3.896
R3943 VSS.n203 VSS.n201 3.896
R3944 VSS.n144 VSS.n142 3.882
R3945 VSS.n147 VSS.n145 3.882
R3946 VSS.n150 VSS.n148 3.882
R3947 VSS.n153 VSS.n151 3.882
R3948 VSS.n156 VSS.n154 3.882
R3949 VSS.n159 VSS.n157 3.882
R3950 VSS.n162 VSS.n160 3.882
R3951 VSS.n165 VSS.n163 3.882
R3952 VSS.n168 VSS.n166 3.882
R3953 VSS.n171 VSS.n169 3.882
R3954 VSS.n174 VSS.n172 3.882
R3955 VSS.n177 VSS.n175 3.882
R3956 VSS.n180 VSS.n178 3.882
R3957 VSS.n183 VSS.n181 3.882
R3958 VSS.n186 VSS.n184 3.882
R3959 VSS.n201 VSS.n194 3.88
R3960 VSS.n142 VSS.n141 3.866
R3961 VSS.n7 VSS.n6 3.827
R3962 VSS.n10 VSS.n4 3.826
R3963 VSS.n2337 VSS.n2336 3.651
R3964 VSS.n1086 VSS.n1085 3.312
R3965 VSS.n1088 VSS.n1087 3.312
R3966 VSS.n1090 VSS.n1089 3.312
R3967 VSS.n1092 VSS.n1091 3.312
R3968 VSS.n1094 VSS.n1093 3.312
R3969 VSS.n1096 VSS.n1095 3.312
R3970 VSS.n1098 VSS.n1097 3.312
R3971 VSS.n1100 VSS.n1099 3.312
R3972 VSS.n1102 VSS.n1101 3.312
R3973 VSS.n1104 VSS.n1103 3.312
R3974 VSS.n1106 VSS.n1105 3.312
R3975 VSS.n1108 VSS.n1107 3.312
R3976 VSS.n1110 VSS.n1109 3.312
R3977 VSS.n1114 VSS.n1111 3.312
R3978 VSS.n1116 VSS.n1115 3.312
R3979 VSS.n1615 VSS.n1614 3.312
R3980 VSS.n1617 VSS.n1616 3.312
R3981 VSS.n1619 VSS.n1618 3.312
R3982 VSS.n1621 VSS.n1620 3.312
R3983 VSS.n1623 VSS.n1622 3.312
R3984 VSS.n1625 VSS.n1624 3.312
R3985 VSS.n1627 VSS.n1626 3.312
R3986 VSS.n1629 VSS.n1628 3.312
R3987 VSS.n1631 VSS.n1630 3.312
R3988 VSS.n1633 VSS.n1632 3.312
R3989 VSS.n1635 VSS.n1634 3.312
R3990 VSS.n1637 VSS.n1636 3.312
R3991 VSS.n1639 VSS.n1638 3.312
R3992 VSS.n1641 VSS.n1640 3.312
R3993 VSS.n1645 VSS.n1642 3.312
R3994 VSS.n2099 VSS.n2098 3.312
R3995 VSS.n2101 VSS.n2100 3.312
R3996 VSS.n2103 VSS.n2102 3.312
R3997 VSS.n2105 VSS.n2104 3.312
R3998 VSS.n2107 VSS.n2106 3.312
R3999 VSS.n2109 VSS.n2108 3.312
R4000 VSS.n2111 VSS.n2110 3.312
R4001 VSS.n2113 VSS.n2112 3.312
R4002 VSS.n2115 VSS.n2114 3.312
R4003 VSS.n2117 VSS.n2116 3.312
R4004 VSS.n2119 VSS.n2118 3.312
R4005 VSS.n2121 VSS.n2120 3.312
R4006 VSS.n2123 VSS.n2122 3.312
R4007 VSS.n2125 VSS.n2124 3.312
R4008 VSS.n2127 VSS.n2126 3.312
R4009 VSS.n623 VSS.n622 3.312
R4010 VSS.n625 VSS.n624 3.312
R4011 VSS.n627 VSS.n626 3.312
R4012 VSS.n629 VSS.n628 3.312
R4013 VSS.n631 VSS.n630 3.312
R4014 VSS.n633 VSS.n632 3.312
R4015 VSS.n635 VSS.n634 3.312
R4016 VSS.n637 VSS.n636 3.312
R4017 VSS.n639 VSS.n638 3.312
R4018 VSS.n641 VSS.n640 3.312
R4019 VSS.n643 VSS.n642 3.312
R4020 VSS.n645 VSS.n644 3.312
R4021 VSS.n647 VSS.n646 3.312
R4022 VSS.n649 VSS.n648 3.312
R4023 VSS.n651 VSS.n650 3.312
R4024 VSS.n2181 VSS.n2180 3.224
R4025 VSS.n2184 VSS.n2183 3.224
R4026 VSS.n2187 VSS.n2186 3.224
R4027 VSS.n2190 VSS.n2189 3.224
R4028 VSS.n2193 VSS.n2192 3.224
R4029 VSS.n2196 VSS.n2195 3.224
R4030 VSS.n2199 VSS.n2198 3.224
R4031 VSS.n2202 VSS.n2201 3.224
R4032 VSS.n2205 VSS.n2204 3.224
R4033 VSS.n2208 VSS.n2207 3.224
R4034 VSS.n2211 VSS.n2210 3.224
R4035 VSS.n2214 VSS.n2213 3.224
R4036 VSS.n2217 VSS.n2216 3.224
R4037 VSS.n2220 VSS.n2219 3.224
R4038 VSS.n2223 VSS.n2222 3.224
R4039 VSS.n1955 VSS.n1954 3.224
R4040 VSS.n1958 VSS.n1957 3.224
R4041 VSS.n1961 VSS.n1960 3.224
R4042 VSS.n1964 VSS.n1963 3.224
R4043 VSS.n1967 VSS.n1966 3.224
R4044 VSS.n1970 VSS.n1969 3.224
R4045 VSS.n1973 VSS.n1972 3.224
R4046 VSS.n1976 VSS.n1975 3.224
R4047 VSS.n1979 VSS.n1978 3.224
R4048 VSS.n1982 VSS.n1981 3.224
R4049 VSS.n1985 VSS.n1984 3.224
R4050 VSS.n1988 VSS.n1987 3.224
R4051 VSS.n1991 VSS.n1990 3.224
R4052 VSS.n1994 VSS.n1993 3.224
R4053 VSS.n1997 VSS.n1996 3.224
R4054 VSS.n1859 VSS.n1858 3.224
R4055 VSS.n1862 VSS.n1861 3.224
R4056 VSS.n1865 VSS.n1864 3.224
R4057 VSS.n1868 VSS.n1867 3.224
R4058 VSS.n1871 VSS.n1870 3.224
R4059 VSS.n1874 VSS.n1873 3.224
R4060 VSS.n1877 VSS.n1876 3.224
R4061 VSS.n1880 VSS.n1879 3.224
R4062 VSS.n1883 VSS.n1882 3.224
R4063 VSS.n1886 VSS.n1885 3.224
R4064 VSS.n1889 VSS.n1888 3.224
R4065 VSS.n1892 VSS.n1891 3.224
R4066 VSS.n1895 VSS.n1894 3.224
R4067 VSS.n1898 VSS.n1897 3.224
R4068 VSS.n1901 VSS.n1900 3.224
R4069 VSS.n1795 VSS.n1794 3.224
R4070 VSS.n1798 VSS.n1797 3.224
R4071 VSS.n1801 VSS.n1800 3.224
R4072 VSS.n1804 VSS.n1803 3.224
R4073 VSS.n1807 VSS.n1806 3.224
R4074 VSS.n1810 VSS.n1809 3.224
R4075 VSS.n1813 VSS.n1812 3.224
R4076 VSS.n1816 VSS.n1815 3.224
R4077 VSS.n1819 VSS.n1818 3.224
R4078 VSS.n1822 VSS.n1821 3.224
R4079 VSS.n1825 VSS.n1824 3.224
R4080 VSS.n1828 VSS.n1827 3.224
R4081 VSS.n1831 VSS.n1830 3.224
R4082 VSS.n1834 VSS.n1833 3.224
R4083 VSS.n1837 VSS.n1836 3.224
R4084 VSS.n1731 VSS.n1730 3.224
R4085 VSS.n1734 VSS.n1733 3.224
R4086 VSS.n1737 VSS.n1736 3.224
R4087 VSS.n1740 VSS.n1739 3.224
R4088 VSS.n1743 VSS.n1742 3.224
R4089 VSS.n1746 VSS.n1745 3.224
R4090 VSS.n1749 VSS.n1748 3.224
R4091 VSS.n1752 VSS.n1751 3.224
R4092 VSS.n1755 VSS.n1754 3.224
R4093 VSS.n1758 VSS.n1757 3.224
R4094 VSS.n1761 VSS.n1760 3.224
R4095 VSS.n1764 VSS.n1763 3.224
R4096 VSS.n1767 VSS.n1766 3.224
R4097 VSS.n1770 VSS.n1769 3.224
R4098 VSS.n1773 VSS.n1772 3.224
R4099 VSS.n1667 VSS.n1666 3.224
R4100 VSS.n1670 VSS.n1669 3.224
R4101 VSS.n1673 VSS.n1672 3.224
R4102 VSS.n1676 VSS.n1675 3.224
R4103 VSS.n1679 VSS.n1678 3.224
R4104 VSS.n1682 VSS.n1681 3.224
R4105 VSS.n1685 VSS.n1684 3.224
R4106 VSS.n1688 VSS.n1687 3.224
R4107 VSS.n1691 VSS.n1690 3.224
R4108 VSS.n1694 VSS.n1693 3.224
R4109 VSS.n1697 VSS.n1696 3.224
R4110 VSS.n1700 VSS.n1699 3.224
R4111 VSS.n1703 VSS.n1702 3.224
R4112 VSS.n1706 VSS.n1705 3.224
R4113 VSS.n1709 VSS.n1708 3.224
R4114 VSS.n1522 VSS.n1521 3.224
R4115 VSS.n1525 VSS.n1524 3.224
R4116 VSS.n1528 VSS.n1527 3.224
R4117 VSS.n1531 VSS.n1530 3.224
R4118 VSS.n1534 VSS.n1533 3.224
R4119 VSS.n1537 VSS.n1536 3.224
R4120 VSS.n1540 VSS.n1539 3.224
R4121 VSS.n1543 VSS.n1542 3.224
R4122 VSS.n1546 VSS.n1545 3.224
R4123 VSS.n1549 VSS.n1548 3.224
R4124 VSS.n1552 VSS.n1551 3.224
R4125 VSS.n1555 VSS.n1554 3.224
R4126 VSS.n1558 VSS.n1557 3.224
R4127 VSS.n1561 VSS.n1560 3.224
R4128 VSS.n1564 VSS.n1563 3.224
R4129 VSS.n1458 VSS.n1457 3.224
R4130 VSS.n1461 VSS.n1460 3.224
R4131 VSS.n1464 VSS.n1463 3.224
R4132 VSS.n1467 VSS.n1466 3.224
R4133 VSS.n1470 VSS.n1469 3.224
R4134 VSS.n1473 VSS.n1472 3.224
R4135 VSS.n1476 VSS.n1475 3.224
R4136 VSS.n1479 VSS.n1478 3.224
R4137 VSS.n1482 VSS.n1481 3.224
R4138 VSS.n1485 VSS.n1484 3.224
R4139 VSS.n1488 VSS.n1487 3.224
R4140 VSS.n1491 VSS.n1490 3.224
R4141 VSS.n1494 VSS.n1493 3.224
R4142 VSS.n1497 VSS.n1496 3.224
R4143 VSS.n1500 VSS.n1499 3.224
R4144 VSS.n1394 VSS.n1393 3.224
R4145 VSS.n1397 VSS.n1396 3.224
R4146 VSS.n1400 VSS.n1399 3.224
R4147 VSS.n1403 VSS.n1402 3.224
R4148 VSS.n1406 VSS.n1405 3.224
R4149 VSS.n1409 VSS.n1408 3.224
R4150 VSS.n1412 VSS.n1411 3.224
R4151 VSS.n1415 VSS.n1414 3.224
R4152 VSS.n1418 VSS.n1417 3.224
R4153 VSS.n1421 VSS.n1420 3.224
R4154 VSS.n1424 VSS.n1423 3.224
R4155 VSS.n1427 VSS.n1426 3.224
R4156 VSS.n1430 VSS.n1429 3.224
R4157 VSS.n1433 VSS.n1432 3.224
R4158 VSS.n1436 VSS.n1435 3.224
R4159 VSS.n1330 VSS.n1329 3.224
R4160 VSS.n1333 VSS.n1332 3.224
R4161 VSS.n1336 VSS.n1335 3.224
R4162 VSS.n1339 VSS.n1338 3.224
R4163 VSS.n1342 VSS.n1341 3.224
R4164 VSS.n1345 VSS.n1344 3.224
R4165 VSS.n1348 VSS.n1347 3.224
R4166 VSS.n1351 VSS.n1350 3.224
R4167 VSS.n1354 VSS.n1353 3.224
R4168 VSS.n1357 VSS.n1356 3.224
R4169 VSS.n1360 VSS.n1359 3.224
R4170 VSS.n1363 VSS.n1362 3.224
R4171 VSS.n1366 VSS.n1365 3.224
R4172 VSS.n1369 VSS.n1368 3.224
R4173 VSS.n1372 VSS.n1371 3.224
R4174 VSS.n1266 VSS.n1265 3.224
R4175 VSS.n1269 VSS.n1268 3.224
R4176 VSS.n1272 VSS.n1271 3.224
R4177 VSS.n1275 VSS.n1274 3.224
R4178 VSS.n1278 VSS.n1277 3.224
R4179 VSS.n1281 VSS.n1280 3.224
R4180 VSS.n1284 VSS.n1283 3.224
R4181 VSS.n1287 VSS.n1286 3.224
R4182 VSS.n1290 VSS.n1289 3.224
R4183 VSS.n1293 VSS.n1292 3.224
R4184 VSS.n1296 VSS.n1295 3.224
R4185 VSS.n1299 VSS.n1298 3.224
R4186 VSS.n1302 VSS.n1301 3.224
R4187 VSS.n1305 VSS.n1304 3.224
R4188 VSS.n1308 VSS.n1307 3.224
R4189 VSS.n1202 VSS.n1201 3.224
R4190 VSS.n1205 VSS.n1204 3.224
R4191 VSS.n1208 VSS.n1207 3.224
R4192 VSS.n1211 VSS.n1210 3.224
R4193 VSS.n1214 VSS.n1213 3.224
R4194 VSS.n1217 VSS.n1216 3.224
R4195 VSS.n1220 VSS.n1219 3.224
R4196 VSS.n1223 VSS.n1222 3.224
R4197 VSS.n1226 VSS.n1225 3.224
R4198 VSS.n1229 VSS.n1228 3.224
R4199 VSS.n1232 VSS.n1231 3.224
R4200 VSS.n1235 VSS.n1234 3.224
R4201 VSS.n1238 VSS.n1237 3.224
R4202 VSS.n1241 VSS.n1240 3.224
R4203 VSS.n1244 VSS.n1243 3.224
R4204 VSS.n1138 VSS.n1137 3.224
R4205 VSS.n1141 VSS.n1140 3.224
R4206 VSS.n1144 VSS.n1143 3.224
R4207 VSS.n1147 VSS.n1146 3.224
R4208 VSS.n1150 VSS.n1149 3.224
R4209 VSS.n1153 VSS.n1152 3.224
R4210 VSS.n1156 VSS.n1155 3.224
R4211 VSS.n1159 VSS.n1158 3.224
R4212 VSS.n1162 VSS.n1161 3.224
R4213 VSS.n1165 VSS.n1164 3.224
R4214 VSS.n1168 VSS.n1167 3.224
R4215 VSS.n1171 VSS.n1170 3.224
R4216 VSS.n1174 VSS.n1173 3.224
R4217 VSS.n1177 VSS.n1176 3.224
R4218 VSS.n1180 VSS.n1179 3.224
R4219 VSS.n993 VSS.n992 3.224
R4220 VSS.n996 VSS.n995 3.224
R4221 VSS.n999 VSS.n998 3.224
R4222 VSS.n1002 VSS.n1001 3.224
R4223 VSS.n1005 VSS.n1004 3.224
R4224 VSS.n1008 VSS.n1007 3.224
R4225 VSS.n1011 VSS.n1010 3.224
R4226 VSS.n1014 VSS.n1013 3.224
R4227 VSS.n1017 VSS.n1016 3.224
R4228 VSS.n1020 VSS.n1019 3.224
R4229 VSS.n1023 VSS.n1022 3.224
R4230 VSS.n1026 VSS.n1025 3.224
R4231 VSS.n1029 VSS.n1028 3.224
R4232 VSS.n1032 VSS.n1031 3.224
R4233 VSS.n1035 VSS.n1034 3.224
R4234 VSS.n929 VSS.n928 3.224
R4235 VSS.n932 VSS.n931 3.224
R4236 VSS.n935 VSS.n934 3.224
R4237 VSS.n938 VSS.n937 3.224
R4238 VSS.n941 VSS.n940 3.224
R4239 VSS.n944 VSS.n943 3.224
R4240 VSS.n947 VSS.n946 3.224
R4241 VSS.n950 VSS.n949 3.224
R4242 VSS.n953 VSS.n952 3.224
R4243 VSS.n956 VSS.n955 3.224
R4244 VSS.n959 VSS.n958 3.224
R4245 VSS.n962 VSS.n961 3.224
R4246 VSS.n965 VSS.n964 3.224
R4247 VSS.n968 VSS.n967 3.224
R4248 VSS.n971 VSS.n970 3.224
R4249 VSS.n865 VSS.n864 3.224
R4250 VSS.n868 VSS.n867 3.224
R4251 VSS.n871 VSS.n870 3.224
R4252 VSS.n874 VSS.n873 3.224
R4253 VSS.n877 VSS.n876 3.224
R4254 VSS.n880 VSS.n879 3.224
R4255 VSS.n883 VSS.n882 3.224
R4256 VSS.n886 VSS.n885 3.224
R4257 VSS.n889 VSS.n888 3.224
R4258 VSS.n892 VSS.n891 3.224
R4259 VSS.n895 VSS.n894 3.224
R4260 VSS.n898 VSS.n897 3.224
R4261 VSS.n901 VSS.n900 3.224
R4262 VSS.n904 VSS.n903 3.224
R4263 VSS.n907 VSS.n906 3.224
R4264 VSS.n801 VSS.n800 3.224
R4265 VSS.n804 VSS.n803 3.224
R4266 VSS.n807 VSS.n806 3.224
R4267 VSS.n810 VSS.n809 3.224
R4268 VSS.n813 VSS.n812 3.224
R4269 VSS.n816 VSS.n815 3.224
R4270 VSS.n819 VSS.n818 3.224
R4271 VSS.n822 VSS.n821 3.224
R4272 VSS.n825 VSS.n824 3.224
R4273 VSS.n828 VSS.n827 3.224
R4274 VSS.n831 VSS.n830 3.224
R4275 VSS.n834 VSS.n833 3.224
R4276 VSS.n837 VSS.n836 3.224
R4277 VSS.n840 VSS.n839 3.224
R4278 VSS.n843 VSS.n842 3.224
R4279 VSS.n705 VSS.n704 3.224
R4280 VSS.n708 VSS.n707 3.224
R4281 VSS.n711 VSS.n710 3.224
R4282 VSS.n714 VSS.n713 3.224
R4283 VSS.n717 VSS.n716 3.224
R4284 VSS.n720 VSS.n719 3.224
R4285 VSS.n723 VSS.n722 3.224
R4286 VSS.n726 VSS.n725 3.224
R4287 VSS.n729 VSS.n728 3.224
R4288 VSS.n732 VSS.n731 3.224
R4289 VSS.n735 VSS.n734 3.224
R4290 VSS.n738 VSS.n737 3.224
R4291 VSS.n741 VSS.n740 3.224
R4292 VSS.n744 VSS.n743 3.224
R4293 VSS.n747 VSS.n746 3.224
R4294 VSS.n496 VSS.n495 3.224
R4295 VSS.n499 VSS.n498 3.224
R4296 VSS.n502 VSS.n501 3.224
R4297 VSS.n505 VSS.n504 3.224
R4298 VSS.n508 VSS.n507 3.224
R4299 VSS.n511 VSS.n510 3.224
R4300 VSS.n514 VSS.n513 3.224
R4301 VSS.n517 VSS.n516 3.224
R4302 VSS.n520 VSS.n519 3.224
R4303 VSS.n523 VSS.n522 3.224
R4304 VSS.n526 VSS.n525 3.224
R4305 VSS.n529 VSS.n528 3.224
R4306 VSS.n532 VSS.n531 3.224
R4307 VSS.n535 VSS.n534 3.224
R4308 VSS.n538 VSS.n537 3.224
R4309 VSS.n191 VSS.n190 3.008
R4310 VSS.n199 VSS.n198 3.008
R4311 VSS.n208 VSS.n207 3.008
R4312 VSS.n217 VSS.n216 3.008
R4313 VSS.n226 VSS.n225 3.008
R4314 VSS.n235 VSS.n234 3.008
R4315 VSS.n244 VSS.n243 3.008
R4316 VSS.n253 VSS.n252 3.008
R4317 VSS.n262 VSS.n261 3.008
R4318 VSS.n271 VSS.n270 3.008
R4319 VSS.n280 VSS.n279 3.008
R4320 VSS.n289 VSS.n288 3.008
R4321 VSS.n298 VSS.n297 3.008
R4322 VSS.n307 VSS.n306 3.008
R4323 VSS.n316 VSS.n315 3.008
R4324 VSS.n325 VSS.n324 3.008
R4325 VSS.n2333 VSS.n2331 2.573
R4326 VSS.n2291 VSS.n2289 2.569
R4327 VSS.n2294 VSS.n2292 2.569
R4328 VSS.n2297 VSS.n2295 2.569
R4329 VSS.n2300 VSS.n2298 2.569
R4330 VSS.n2303 VSS.n2301 2.569
R4331 VSS.n2306 VSS.n2304 2.569
R4332 VSS.n2309 VSS.n2307 2.569
R4333 VSS.n2312 VSS.n2310 2.569
R4334 VSS.n2315 VSS.n2313 2.569
R4335 VSS.n2318 VSS.n2316 2.569
R4336 VSS.n2321 VSS.n2319 2.569
R4337 VSS.n2324 VSS.n2322 2.569
R4338 VSS.n2327 VSS.n2325 2.569
R4339 VSS.n2330 VSS.n2328 2.569
R4340 VSS.n2334 VSS.n2333 2.316
R4341 VSS.n2292 VSS.n2291 2.313
R4342 VSS.n2295 VSS.n2294 2.313
R4343 VSS.n2298 VSS.n2297 2.313
R4344 VSS.n2301 VSS.n2300 2.313
R4345 VSS.n2304 VSS.n2303 2.313
R4346 VSS.n2307 VSS.n2306 2.313
R4347 VSS.n2310 VSS.n2309 2.313
R4348 VSS.n2313 VSS.n2312 2.313
R4349 VSS.n2316 VSS.n2315 2.313
R4350 VSS.n2319 VSS.n2318 2.313
R4351 VSS.n2322 VSS.n2321 2.313
R4352 VSS.n2325 VSS.n2324 2.313
R4353 VSS.n2328 VSS.n2327 2.313
R4354 VSS.n2331 VSS.n2330 2.313
R4355 VSS.n1710 VSS.n1646 2.235
R4356 VSS.n1181 VSS.n1117 2.227
R4357 VSS.n908 VSS.n844 1.893
R4358 VSS.n972 VSS.n908 1.893
R4359 VSS.n1036 VSS.n972 1.893
R4360 VSS.n1117 VSS.n1036 1.893
R4361 VSS.n1245 VSS.n1181 1.893
R4362 VSS.n1309 VSS.n1245 1.893
R4363 VSS.n1373 VSS.n1309 1.893
R4364 VSS.n1437 VSS.n1373 1.893
R4365 VSS.n1501 VSS.n1437 1.893
R4366 VSS.n1565 VSS.n1501 1.893
R4367 VSS.n1646 VSS.n1565 1.893
R4368 VSS.n1774 VSS.n1710 1.893
R4369 VSS.n1838 VSS.n1774 1.893
R4370 VSS.n1902 VSS.n1838 1.879
R4371 VSS.n1085 VSS.n1084 1.821
R4372 VSS.n1087 VSS.n1086 1.821
R4373 VSS.n1089 VSS.n1088 1.821
R4374 VSS.n1091 VSS.n1090 1.821
R4375 VSS.n1093 VSS.n1092 1.821
R4376 VSS.n1095 VSS.n1094 1.821
R4377 VSS.n1097 VSS.n1096 1.821
R4378 VSS.n1099 VSS.n1098 1.821
R4379 VSS.n1101 VSS.n1100 1.821
R4380 VSS.n1103 VSS.n1102 1.821
R4381 VSS.n1105 VSS.n1104 1.821
R4382 VSS.n1107 VSS.n1106 1.821
R4383 VSS.n1109 VSS.n1108 1.821
R4384 VSS.n1111 VSS.n1110 1.821
R4385 VSS.n1115 VSS.n1114 1.821
R4386 VSS.n1614 VSS.n1613 1.821
R4387 VSS.n1616 VSS.n1615 1.821
R4388 VSS.n1618 VSS.n1617 1.821
R4389 VSS.n1620 VSS.n1619 1.821
R4390 VSS.n1622 VSS.n1621 1.821
R4391 VSS.n1624 VSS.n1623 1.821
R4392 VSS.n1626 VSS.n1625 1.821
R4393 VSS.n1628 VSS.n1627 1.821
R4394 VSS.n1630 VSS.n1629 1.821
R4395 VSS.n1632 VSS.n1631 1.821
R4396 VSS.n1634 VSS.n1633 1.821
R4397 VSS.n1636 VSS.n1635 1.821
R4398 VSS.n1638 VSS.n1637 1.821
R4399 VSS.n1640 VSS.n1639 1.821
R4400 VSS.n1642 VSS.n1641 1.821
R4401 VSS.n2098 VSS.n2097 1.821
R4402 VSS.n2100 VSS.n2099 1.821
R4403 VSS.n2102 VSS.n2101 1.821
R4404 VSS.n2104 VSS.n2103 1.821
R4405 VSS.n2106 VSS.n2105 1.821
R4406 VSS.n2108 VSS.n2107 1.821
R4407 VSS.n2110 VSS.n2109 1.821
R4408 VSS.n2112 VSS.n2111 1.821
R4409 VSS.n2114 VSS.n2113 1.821
R4410 VSS.n2116 VSS.n2115 1.821
R4411 VSS.n2118 VSS.n2117 1.821
R4412 VSS.n2120 VSS.n2119 1.821
R4413 VSS.n2122 VSS.n2121 1.821
R4414 VSS.n2124 VSS.n2123 1.821
R4415 VSS.n2126 VSS.n2125 1.821
R4416 VSS.n622 VSS.n621 1.821
R4417 VSS.n624 VSS.n623 1.821
R4418 VSS.n626 VSS.n625 1.821
R4419 VSS.n628 VSS.n627 1.821
R4420 VSS.n630 VSS.n629 1.821
R4421 VSS.n632 VSS.n631 1.821
R4422 VSS.n634 VSS.n633 1.821
R4423 VSS.n636 VSS.n635 1.821
R4424 VSS.n638 VSS.n637 1.821
R4425 VSS.n640 VSS.n639 1.821
R4426 VSS.n642 VSS.n641 1.821
R4427 VSS.n644 VSS.n643 1.821
R4428 VSS.n646 VSS.n645 1.821
R4429 VSS.n648 VSS.n647 1.821
R4430 VSS.n650 VSS.n649 1.821
R4431 VSS.n345 VSS.n344 1.816
R4432 VSS.n347 VSS.n346 1.798
R4433 VSS.n349 VSS.n348 1.786
R4434 VSS.n344 VSS.n343 1.78
R4435 VSS.n348 VSS.n347 1.776
R4436 VSS.n346 VSS.n345 1.772
R4437 VSS.n2180 VSS.n2178 1.745
R4438 VSS.n2183 VSS.n2181 1.745
R4439 VSS.n2186 VSS.n2184 1.745
R4440 VSS.n2189 VSS.n2187 1.745
R4441 VSS.n2192 VSS.n2190 1.745
R4442 VSS.n2195 VSS.n2193 1.745
R4443 VSS.n2198 VSS.n2196 1.745
R4444 VSS.n2201 VSS.n2199 1.745
R4445 VSS.n2204 VSS.n2202 1.745
R4446 VSS.n2207 VSS.n2205 1.745
R4447 VSS.n2210 VSS.n2208 1.745
R4448 VSS.n2213 VSS.n2211 1.745
R4449 VSS.n2216 VSS.n2214 1.745
R4450 VSS.n2219 VSS.n2217 1.745
R4451 VSS.n2222 VSS.n2220 1.745
R4452 VSS.n1954 VSS.n1952 1.745
R4453 VSS.n1957 VSS.n1955 1.745
R4454 VSS.n1960 VSS.n1958 1.745
R4455 VSS.n1963 VSS.n1961 1.745
R4456 VSS.n1966 VSS.n1964 1.745
R4457 VSS.n1969 VSS.n1967 1.745
R4458 VSS.n1972 VSS.n1970 1.745
R4459 VSS.n1975 VSS.n1973 1.745
R4460 VSS.n1978 VSS.n1976 1.745
R4461 VSS.n1981 VSS.n1979 1.745
R4462 VSS.n1984 VSS.n1982 1.745
R4463 VSS.n1987 VSS.n1985 1.745
R4464 VSS.n1990 VSS.n1988 1.745
R4465 VSS.n1993 VSS.n1991 1.745
R4466 VSS.n1996 VSS.n1994 1.745
R4467 VSS.n1858 VSS.n1856 1.745
R4468 VSS.n1861 VSS.n1859 1.745
R4469 VSS.n1864 VSS.n1862 1.745
R4470 VSS.n1867 VSS.n1865 1.745
R4471 VSS.n1870 VSS.n1868 1.745
R4472 VSS.n1873 VSS.n1871 1.745
R4473 VSS.n1876 VSS.n1874 1.745
R4474 VSS.n1879 VSS.n1877 1.745
R4475 VSS.n1882 VSS.n1880 1.745
R4476 VSS.n1885 VSS.n1883 1.745
R4477 VSS.n1888 VSS.n1886 1.745
R4478 VSS.n1891 VSS.n1889 1.745
R4479 VSS.n1894 VSS.n1892 1.745
R4480 VSS.n1897 VSS.n1895 1.745
R4481 VSS.n1900 VSS.n1898 1.745
R4482 VSS.n1794 VSS.n1792 1.745
R4483 VSS.n1797 VSS.n1795 1.745
R4484 VSS.n1800 VSS.n1798 1.745
R4485 VSS.n1803 VSS.n1801 1.745
R4486 VSS.n1806 VSS.n1804 1.745
R4487 VSS.n1809 VSS.n1807 1.745
R4488 VSS.n1812 VSS.n1810 1.745
R4489 VSS.n1815 VSS.n1813 1.745
R4490 VSS.n1818 VSS.n1816 1.745
R4491 VSS.n1821 VSS.n1819 1.745
R4492 VSS.n1824 VSS.n1822 1.745
R4493 VSS.n1827 VSS.n1825 1.745
R4494 VSS.n1830 VSS.n1828 1.745
R4495 VSS.n1833 VSS.n1831 1.745
R4496 VSS.n1836 VSS.n1834 1.745
R4497 VSS.n1730 VSS.n1728 1.745
R4498 VSS.n1733 VSS.n1731 1.745
R4499 VSS.n1736 VSS.n1734 1.745
R4500 VSS.n1739 VSS.n1737 1.745
R4501 VSS.n1742 VSS.n1740 1.745
R4502 VSS.n1745 VSS.n1743 1.745
R4503 VSS.n1748 VSS.n1746 1.745
R4504 VSS.n1751 VSS.n1749 1.745
R4505 VSS.n1754 VSS.n1752 1.745
R4506 VSS.n1757 VSS.n1755 1.745
R4507 VSS.n1760 VSS.n1758 1.745
R4508 VSS.n1763 VSS.n1761 1.745
R4509 VSS.n1766 VSS.n1764 1.745
R4510 VSS.n1769 VSS.n1767 1.745
R4511 VSS.n1772 VSS.n1770 1.745
R4512 VSS.n1666 VSS.n1664 1.745
R4513 VSS.n1669 VSS.n1667 1.745
R4514 VSS.n1672 VSS.n1670 1.745
R4515 VSS.n1675 VSS.n1673 1.745
R4516 VSS.n1678 VSS.n1676 1.745
R4517 VSS.n1681 VSS.n1679 1.745
R4518 VSS.n1684 VSS.n1682 1.745
R4519 VSS.n1687 VSS.n1685 1.745
R4520 VSS.n1690 VSS.n1688 1.745
R4521 VSS.n1693 VSS.n1691 1.745
R4522 VSS.n1696 VSS.n1694 1.745
R4523 VSS.n1699 VSS.n1697 1.745
R4524 VSS.n1702 VSS.n1700 1.745
R4525 VSS.n1705 VSS.n1703 1.745
R4526 VSS.n1708 VSS.n1706 1.745
R4527 VSS.n1521 VSS.n1519 1.745
R4528 VSS.n1524 VSS.n1522 1.745
R4529 VSS.n1527 VSS.n1525 1.745
R4530 VSS.n1530 VSS.n1528 1.745
R4531 VSS.n1533 VSS.n1531 1.745
R4532 VSS.n1536 VSS.n1534 1.745
R4533 VSS.n1539 VSS.n1537 1.745
R4534 VSS.n1542 VSS.n1540 1.745
R4535 VSS.n1545 VSS.n1543 1.745
R4536 VSS.n1548 VSS.n1546 1.745
R4537 VSS.n1551 VSS.n1549 1.745
R4538 VSS.n1554 VSS.n1552 1.745
R4539 VSS.n1557 VSS.n1555 1.745
R4540 VSS.n1560 VSS.n1558 1.745
R4541 VSS.n1563 VSS.n1561 1.745
R4542 VSS.n1457 VSS.n1455 1.745
R4543 VSS.n1460 VSS.n1458 1.745
R4544 VSS.n1463 VSS.n1461 1.745
R4545 VSS.n1466 VSS.n1464 1.745
R4546 VSS.n1469 VSS.n1467 1.745
R4547 VSS.n1472 VSS.n1470 1.745
R4548 VSS.n1475 VSS.n1473 1.745
R4549 VSS.n1478 VSS.n1476 1.745
R4550 VSS.n1481 VSS.n1479 1.745
R4551 VSS.n1484 VSS.n1482 1.745
R4552 VSS.n1487 VSS.n1485 1.745
R4553 VSS.n1490 VSS.n1488 1.745
R4554 VSS.n1493 VSS.n1491 1.745
R4555 VSS.n1496 VSS.n1494 1.745
R4556 VSS.n1499 VSS.n1497 1.745
R4557 VSS.n1393 VSS.n1391 1.745
R4558 VSS.n1396 VSS.n1394 1.745
R4559 VSS.n1399 VSS.n1397 1.745
R4560 VSS.n1402 VSS.n1400 1.745
R4561 VSS.n1405 VSS.n1403 1.745
R4562 VSS.n1408 VSS.n1406 1.745
R4563 VSS.n1411 VSS.n1409 1.745
R4564 VSS.n1414 VSS.n1412 1.745
R4565 VSS.n1417 VSS.n1415 1.745
R4566 VSS.n1420 VSS.n1418 1.745
R4567 VSS.n1423 VSS.n1421 1.745
R4568 VSS.n1426 VSS.n1424 1.745
R4569 VSS.n1429 VSS.n1427 1.745
R4570 VSS.n1432 VSS.n1430 1.745
R4571 VSS.n1435 VSS.n1433 1.745
R4572 VSS.n1329 VSS.n1327 1.745
R4573 VSS.n1332 VSS.n1330 1.745
R4574 VSS.n1335 VSS.n1333 1.745
R4575 VSS.n1338 VSS.n1336 1.745
R4576 VSS.n1341 VSS.n1339 1.745
R4577 VSS.n1344 VSS.n1342 1.745
R4578 VSS.n1347 VSS.n1345 1.745
R4579 VSS.n1350 VSS.n1348 1.745
R4580 VSS.n1353 VSS.n1351 1.745
R4581 VSS.n1356 VSS.n1354 1.745
R4582 VSS.n1359 VSS.n1357 1.745
R4583 VSS.n1362 VSS.n1360 1.745
R4584 VSS.n1365 VSS.n1363 1.745
R4585 VSS.n1368 VSS.n1366 1.745
R4586 VSS.n1371 VSS.n1369 1.745
R4587 VSS.n1265 VSS.n1263 1.745
R4588 VSS.n1268 VSS.n1266 1.745
R4589 VSS.n1271 VSS.n1269 1.745
R4590 VSS.n1274 VSS.n1272 1.745
R4591 VSS.n1277 VSS.n1275 1.745
R4592 VSS.n1280 VSS.n1278 1.745
R4593 VSS.n1283 VSS.n1281 1.745
R4594 VSS.n1286 VSS.n1284 1.745
R4595 VSS.n1289 VSS.n1287 1.745
R4596 VSS.n1292 VSS.n1290 1.745
R4597 VSS.n1295 VSS.n1293 1.745
R4598 VSS.n1298 VSS.n1296 1.745
R4599 VSS.n1301 VSS.n1299 1.745
R4600 VSS.n1304 VSS.n1302 1.745
R4601 VSS.n1307 VSS.n1305 1.745
R4602 VSS.n1201 VSS.n1199 1.745
R4603 VSS.n1204 VSS.n1202 1.745
R4604 VSS.n1207 VSS.n1205 1.745
R4605 VSS.n1210 VSS.n1208 1.745
R4606 VSS.n1213 VSS.n1211 1.745
R4607 VSS.n1216 VSS.n1214 1.745
R4608 VSS.n1219 VSS.n1217 1.745
R4609 VSS.n1222 VSS.n1220 1.745
R4610 VSS.n1225 VSS.n1223 1.745
R4611 VSS.n1228 VSS.n1226 1.745
R4612 VSS.n1231 VSS.n1229 1.745
R4613 VSS.n1234 VSS.n1232 1.745
R4614 VSS.n1237 VSS.n1235 1.745
R4615 VSS.n1240 VSS.n1238 1.745
R4616 VSS.n1243 VSS.n1241 1.745
R4617 VSS.n1137 VSS.n1135 1.745
R4618 VSS.n1140 VSS.n1138 1.745
R4619 VSS.n1143 VSS.n1141 1.745
R4620 VSS.n1146 VSS.n1144 1.745
R4621 VSS.n1149 VSS.n1147 1.745
R4622 VSS.n1152 VSS.n1150 1.745
R4623 VSS.n1155 VSS.n1153 1.745
R4624 VSS.n1158 VSS.n1156 1.745
R4625 VSS.n1161 VSS.n1159 1.745
R4626 VSS.n1164 VSS.n1162 1.745
R4627 VSS.n1167 VSS.n1165 1.745
R4628 VSS.n1170 VSS.n1168 1.745
R4629 VSS.n1173 VSS.n1171 1.745
R4630 VSS.n1176 VSS.n1174 1.745
R4631 VSS.n1179 VSS.n1177 1.745
R4632 VSS.n992 VSS.n990 1.745
R4633 VSS.n995 VSS.n993 1.745
R4634 VSS.n998 VSS.n996 1.745
R4635 VSS.n1001 VSS.n999 1.745
R4636 VSS.n1004 VSS.n1002 1.745
R4637 VSS.n1007 VSS.n1005 1.745
R4638 VSS.n1010 VSS.n1008 1.745
R4639 VSS.n1013 VSS.n1011 1.745
R4640 VSS.n1016 VSS.n1014 1.745
R4641 VSS.n1019 VSS.n1017 1.745
R4642 VSS.n1022 VSS.n1020 1.745
R4643 VSS.n1025 VSS.n1023 1.745
R4644 VSS.n1028 VSS.n1026 1.745
R4645 VSS.n1031 VSS.n1029 1.745
R4646 VSS.n1034 VSS.n1032 1.745
R4647 VSS.n928 VSS.n926 1.745
R4648 VSS.n931 VSS.n929 1.745
R4649 VSS.n934 VSS.n932 1.745
R4650 VSS.n937 VSS.n935 1.745
R4651 VSS.n940 VSS.n938 1.745
R4652 VSS.n943 VSS.n941 1.745
R4653 VSS.n946 VSS.n944 1.745
R4654 VSS.n949 VSS.n947 1.745
R4655 VSS.n952 VSS.n950 1.745
R4656 VSS.n955 VSS.n953 1.745
R4657 VSS.n958 VSS.n956 1.745
R4658 VSS.n961 VSS.n959 1.745
R4659 VSS.n964 VSS.n962 1.745
R4660 VSS.n967 VSS.n965 1.745
R4661 VSS.n970 VSS.n968 1.745
R4662 VSS.n864 VSS.n862 1.745
R4663 VSS.n867 VSS.n865 1.745
R4664 VSS.n870 VSS.n868 1.745
R4665 VSS.n873 VSS.n871 1.745
R4666 VSS.n876 VSS.n874 1.745
R4667 VSS.n879 VSS.n877 1.745
R4668 VSS.n882 VSS.n880 1.745
R4669 VSS.n885 VSS.n883 1.745
R4670 VSS.n888 VSS.n886 1.745
R4671 VSS.n891 VSS.n889 1.745
R4672 VSS.n894 VSS.n892 1.745
R4673 VSS.n897 VSS.n895 1.745
R4674 VSS.n900 VSS.n898 1.745
R4675 VSS.n903 VSS.n901 1.745
R4676 VSS.n906 VSS.n904 1.745
R4677 VSS.n800 VSS.n798 1.745
R4678 VSS.n803 VSS.n801 1.745
R4679 VSS.n806 VSS.n804 1.745
R4680 VSS.n809 VSS.n807 1.745
R4681 VSS.n812 VSS.n810 1.745
R4682 VSS.n815 VSS.n813 1.745
R4683 VSS.n818 VSS.n816 1.745
R4684 VSS.n821 VSS.n819 1.745
R4685 VSS.n824 VSS.n822 1.745
R4686 VSS.n827 VSS.n825 1.745
R4687 VSS.n830 VSS.n828 1.745
R4688 VSS.n833 VSS.n831 1.745
R4689 VSS.n836 VSS.n834 1.745
R4690 VSS.n839 VSS.n837 1.745
R4691 VSS.n842 VSS.n840 1.745
R4692 VSS.n704 VSS.n702 1.745
R4693 VSS.n707 VSS.n705 1.745
R4694 VSS.n710 VSS.n708 1.745
R4695 VSS.n713 VSS.n711 1.745
R4696 VSS.n716 VSS.n714 1.745
R4697 VSS.n719 VSS.n717 1.745
R4698 VSS.n722 VSS.n720 1.745
R4699 VSS.n725 VSS.n723 1.745
R4700 VSS.n728 VSS.n726 1.745
R4701 VSS.n731 VSS.n729 1.745
R4702 VSS.n734 VSS.n732 1.745
R4703 VSS.n737 VSS.n735 1.745
R4704 VSS.n740 VSS.n738 1.745
R4705 VSS.n743 VSS.n741 1.745
R4706 VSS.n746 VSS.n744 1.745
R4707 VSS.n495 VSS.n493 1.745
R4708 VSS.n498 VSS.n496 1.745
R4709 VSS.n501 VSS.n499 1.745
R4710 VSS.n504 VSS.n502 1.745
R4711 VSS.n507 VSS.n505 1.745
R4712 VSS.n510 VSS.n508 1.745
R4713 VSS.n513 VSS.n511 1.745
R4714 VSS.n516 VSS.n514 1.745
R4715 VSS.n519 VSS.n517 1.745
R4716 VSS.n522 VSS.n520 1.745
R4717 VSS.n525 VSS.n523 1.745
R4718 VSS.n528 VSS.n526 1.745
R4719 VSS.n531 VSS.n529 1.745
R4720 VSS.n534 VSS.n532 1.745
R4721 VSS.n537 VSS.n535 1.745
R4722 VSS.n2337 VSS.n349 1.719
R4723 VSS.n352 VSS.n351 1.552
R4724 VSS.n354 VSS.n353 1.552
R4725 VSS.n356 VSS.n355 1.552
R4726 VSS.n358 VSS.n357 1.552
R4727 VSS.n360 VSS.n359 1.552
R4728 VSS.n362 VSS.n361 1.552
R4729 VSS.n364 VSS.n363 1.552
R4730 VSS.n366 VSS.n365 1.552
R4731 VSS.n368 VSS.n367 1.552
R4732 VSS.n370 VSS.n369 1.552
R4733 VSS.n372 VSS.n371 1.552
R4734 VSS.n374 VSS.n373 1.552
R4735 VSS.n376 VSS.n375 1.552
R4736 VSS.n378 VSS.n377 1.552
R4737 VSS.n380 VSS.n379 1.552
R4738 VSS.n382 VSS.n381 1.552
R4739 VSS.n384 VSS.n383 1.552
R4740 VSS.n386 VSS.n385 1.552
R4741 VSS.n388 VSS.n387 1.552
R4742 VSS.n390 VSS.n389 1.552
R4743 VSS.n392 VSS.n391 1.552
R4744 VSS.n394 VSS.n393 1.552
R4745 VSS.n396 VSS.n395 1.552
R4746 VSS.n398 VSS.n397 1.552
R4747 VSS.n400 VSS.n399 1.552
R4748 VSS.n402 VSS.n401 1.552
R4749 VSS.n404 VSS.n403 1.552
R4750 VSS.n406 VSS.n405 1.552
R4751 VSS.n408 VSS.n407 1.552
R4752 VSS.n410 VSS.n409 1.552
R4753 VSS.n412 VSS.n411 1.552
R4754 VSS.n2336 VSS.n412 1.461
R4755 VSS.n334 VSS.n139 1.335
R4756 VSS.n353 VSS.n352 1.178
R4757 VSS.n357 VSS.n356 1.178
R4758 VSS.n361 VSS.n360 1.178
R4759 VSS.n365 VSS.n364 1.178
R4760 VSS.n369 VSS.n368 1.178
R4761 VSS.n373 VSS.n372 1.178
R4762 VSS.n377 VSS.n376 1.178
R4763 VSS.n381 VSS.n380 1.178
R4764 VSS.n385 VSS.n384 1.178
R4765 VSS.n389 VSS.n388 1.178
R4766 VSS.n393 VSS.n392 1.178
R4767 VSS.n397 VSS.n396 1.178
R4768 VSS.n401 VSS.n400 1.178
R4769 VSS.n405 VSS.n404 1.178
R4770 VSS.n409 VSS.n408 1.178
R4771 VSS.n2144 VSS.n2128 1.063
R4772 VSS.n668 VSS.n652 1.013
R4773 VSS.n2091 VSS.t34 0.732
R4774 VSS.n2087 VSS.t51 0.732
R4775 VSS.n2083 VSS.t35 0.732
R4776 VSS.n2079 VSS.t53 0.732
R4777 VSS.n2075 VSS.t52 0.732
R4778 VSS.n2071 VSS.t4 0.732
R4779 VSS.n2067 VSS.t33 0.732
R4780 VSS.n2063 VSS.t32 0.732
R4781 VSS.n2059 VSS.t5 0.732
R4782 VSS.n2055 VSS.t37 0.732
R4783 VSS.n2051 VSS.t43 0.732
R4784 VSS.n2047 VSS.t31 0.732
R4785 VSS.n2043 VSS.t86 0.732
R4786 VSS.n2039 VSS.t36 0.732
R4787 VSS.n2035 VSS.t42 0.732
R4788 VSS.n2031 VSS.t38 0.732
R4789 VSS.n2256 VSS.n2240 0.582
R4790 VSS VSS.n2338 0.582
R4791 VSS.n555 VSS.n539 0.579
R4792 VSS.n475 VSS.n459 0.574
R4793 VSS.n684 VSS.n668 0.574
R4794 VSS.n1918 VSS.n1902 0.565
R4795 VSS.n764 VSS.n748 0.563
R4796 VSS.n780 VSS.n764 0.557
R4797 VSS.n2014 VSS.n1998 0.553
R4798 VSS.n2128 VSS.n2030 0.538
R4799 VSS.n571 VSS.n555 0.524
R4800 VSS.n2160 VSS.n2144 0.524
R4801 VSS.n2240 VSS.n2224 0.524
R4802 VSS.n1934 VSS.n1918 0.515
R4803 VSS.n2030 VSS.n2014 0.515
R4804 VSS.n1998 VSS.n1934 0.512
R4805 VSS.n652 VSS.n571 0.504
R4806 VSS.n2224 VSS.n2160 0.499
R4807 VSS.n748 VSS.n684 0.488
R4808 VSS.n844 VSS.n780 0.488
R4809 VSS.n2288 VSS.n2256 0.488
R4810 VSS.n539 VSS.n475 0.471
R4811 VSS.n351 VSS.n350 0.348
R4812 VSS.n355 VSS.n354 0.348
R4813 VSS.n359 VSS.n358 0.348
R4814 VSS.n363 VSS.n362 0.348
R4815 VSS.n367 VSS.n366 0.348
R4816 VSS.n371 VSS.n370 0.348
R4817 VSS.n375 VSS.n374 0.348
R4818 VSS.n379 VSS.n378 0.348
R4819 VSS.n383 VSS.n382 0.348
R4820 VSS.n387 VSS.n386 0.348
R4821 VSS.n391 VSS.n390 0.348
R4822 VSS.n395 VSS.n394 0.348
R4823 VSS.n399 VSS.n398 0.348
R4824 VSS.n403 VSS.n402 0.348
R4825 VSS.n407 VSS.n406 0.348
R4826 VSS.n411 VSS.n410 0.348
R4827 VSS.n200 VSS.n199 0.048
R4828 VSS.n209 VSS.n208 0.048
R4829 VSS.n218 VSS.n217 0.048
R4830 VSS.n227 VSS.n226 0.048
R4831 VSS.n236 VSS.n235 0.048
R4832 VSS.n245 VSS.n244 0.048
R4833 VSS.n254 VSS.n253 0.048
R4834 VSS.n263 VSS.n262 0.048
R4835 VSS.n272 VSS.n271 0.048
R4836 VSS.n281 VSS.n280 0.048
R4837 VSS.n290 VSS.n289 0.048
R4838 VSS.n299 VSS.n298 0.048
R4839 VSS.n308 VSS.n307 0.048
R4840 VSS.n317 VSS.n316 0.048
R4841 VSS.n326 VSS.n325 0.048
R4842 VSS.n192 VSS.n191 0.048
R4843 VSS.n199 VSS.n195 0.028
R4844 VSS.n208 VSS.n204 0.028
R4845 VSS.n217 VSS.n213 0.028
R4846 VSS.n226 VSS.n222 0.028
R4847 VSS.n235 VSS.n231 0.028
R4848 VSS.n244 VSS.n240 0.028
R4849 VSS.n253 VSS.n249 0.028
R4850 VSS.n262 VSS.n258 0.028
R4851 VSS.n271 VSS.n267 0.028
R4852 VSS.n280 VSS.n276 0.028
R4853 VSS.n289 VSS.n285 0.028
R4854 VSS.n298 VSS.n294 0.028
R4855 VSS.n307 VSS.n303 0.028
R4856 VSS.n316 VSS.n312 0.028
R4857 VSS.n325 VSS.n321 0.028
R4858 VSS.n191 VSS.n187 0.028
R4859 VSS.n190 VSS.n188 0.003
R4860 VSS.n198 VSS.n196 0.003
R4861 VSS.n207 VSS.n205 0.003
R4862 VSS.n216 VSS.n214 0.003
R4863 VSS.n225 VSS.n223 0.003
R4864 VSS.n234 VSS.n232 0.003
R4865 VSS.n243 VSS.n241 0.003
R4866 VSS.n252 VSS.n250 0.003
R4867 VSS.n261 VSS.n259 0.003
R4868 VSS.n270 VSS.n268 0.003
R4869 VSS.n279 VSS.n277 0.003
R4870 VSS.n288 VSS.n286 0.003
R4871 VSS.n297 VSS.n295 0.003
R4872 VSS.n306 VSS.n304 0.003
R4873 VSS.n315 VSS.n313 0.003
R4874 VSS.n324 VSS.n322 0.003
R4875 a_2015_2180.t0 a_2015_2180.t1 242.857
R4876 PRE_VLSA.n154 PRE_VLSA.t35 572.725
R4877 PRE_VLSA.n144 PRE_VLSA.t22 572.725
R4878 PRE_VLSA.n134 PRE_VLSA.t32 572.725
R4879 PRE_VLSA.n124 PRE_VLSA.t10 572.725
R4880 PRE_VLSA.n114 PRE_VLSA.t14 572.725
R4881 PRE_VLSA.n104 PRE_VLSA.t42 572.725
R4882 PRE_VLSA.n94 PRE_VLSA.t15 572.725
R4883 PRE_VLSA.n84 PRE_VLSA.t44 572.725
R4884 PRE_VLSA.n74 PRE_VLSA.t47 572.725
R4885 PRE_VLSA.n64 PRE_VLSA.t27 572.725
R4886 PRE_VLSA.n54 PRE_VLSA.t43 572.725
R4887 PRE_VLSA.n44 PRE_VLSA.t29 572.725
R4888 PRE_VLSA.n34 PRE_VLSA.t26 572.725
R4889 PRE_VLSA.n24 PRE_VLSA.t11 572.725
R4890 PRE_VLSA.n14 PRE_VLSA.t28 572.725
R4891 PRE_VLSA.n4 PRE_VLSA.t8 572.725
R4892 PRE_VLSA.n0 PRE_VLSA.t13 536.375
R4893 PRE_VLSA.n8 PRE_VLSA.t38 534.877
R4894 PRE_VLSA.n18 PRE_VLSA.t12 534.877
R4895 PRE_VLSA.n28 PRE_VLSA.t5 534.877
R4896 PRE_VLSA.n38 PRE_VLSA.t30 534.877
R4897 PRE_VLSA.n48 PRE_VLSA.t2 534.877
R4898 PRE_VLSA.n58 PRE_VLSA.t36 534.877
R4899 PRE_VLSA.n68 PRE_VLSA.t19 534.877
R4900 PRE_VLSA.n78 PRE_VLSA.t3 534.877
R4901 PRE_VLSA.n88 PRE_VLSA.t17 534.877
R4902 PRE_VLSA.n98 PRE_VLSA.t0 534.877
R4903 PRE_VLSA.n108 PRE_VLSA.t33 534.877
R4904 PRE_VLSA.n118 PRE_VLSA.t18 534.877
R4905 PRE_VLSA.n128 PRE_VLSA.t41 534.877
R4906 PRE_VLSA.n138 PRE_VLSA.t16 534.877
R4907 PRE_VLSA.n148 PRE_VLSA.t9 534.877
R4908 PRE_VLSA.n153 PRE_VLSA.t7 534.866
R4909 PRE_VLSA.n3 PRE_VLSA.t6 534.866
R4910 PRE_VLSA.n13 PRE_VLSA.t31 534.866
R4911 PRE_VLSA.n23 PRE_VLSA.t24 534.866
R4912 PRE_VLSA.n33 PRE_VLSA.t46 534.866
R4913 PRE_VLSA.n43 PRE_VLSA.t21 534.866
R4914 PRE_VLSA.n53 PRE_VLSA.t45 534.866
R4915 PRE_VLSA.n63 PRE_VLSA.t40 534.866
R4916 PRE_VLSA.n73 PRE_VLSA.t23 534.866
R4917 PRE_VLSA.n83 PRE_VLSA.t37 534.866
R4918 PRE_VLSA.n93 PRE_VLSA.t20 534.866
R4919 PRE_VLSA.n103 PRE_VLSA.t4 534.866
R4920 PRE_VLSA.n113 PRE_VLSA.t39 534.866
R4921 PRE_VLSA.n123 PRE_VLSA.t1 534.866
R4922 PRE_VLSA.n133 PRE_VLSA.t34 534.866
R4923 PRE_VLSA.n143 PRE_VLSA.t25 534.866
R4924 PRE_VLSA PRE_VLSA.n155 43.625
R4925 PRE_VLSA.n1 PRE_VLSA.n0 3.102
R4926 PRE_VLSA.n11 PRE_VLSA.n10 3.067
R4927 PRE_VLSA.n21 PRE_VLSA.n20 3.067
R4928 PRE_VLSA.n31 PRE_VLSA.n30 3.067
R4929 PRE_VLSA.n41 PRE_VLSA.n40 3.067
R4930 PRE_VLSA.n51 PRE_VLSA.n50 3.067
R4931 PRE_VLSA.n61 PRE_VLSA.n60 3.067
R4932 PRE_VLSA.n71 PRE_VLSA.n70 3.067
R4933 PRE_VLSA.n81 PRE_VLSA.n80 3.067
R4934 PRE_VLSA.n91 PRE_VLSA.n90 3.067
R4935 PRE_VLSA.n101 PRE_VLSA.n100 3.067
R4936 PRE_VLSA.n111 PRE_VLSA.n110 3.067
R4937 PRE_VLSA.n121 PRE_VLSA.n120 3.067
R4938 PRE_VLSA.n131 PRE_VLSA.n130 3.067
R4939 PRE_VLSA.n141 PRE_VLSA.n140 3.067
R4940 PRE_VLSA.n151 PRE_VLSA.n150 3.046
R4941 PRE_VLSA.n4 PRE_VLSA.n3 2.992
R4942 PRE_VLSA.n9 PRE_VLSA.n8 2.992
R4943 PRE_VLSA.n14 PRE_VLSA.n13 2.992
R4944 PRE_VLSA.n19 PRE_VLSA.n18 2.992
R4945 PRE_VLSA.n24 PRE_VLSA.n23 2.992
R4946 PRE_VLSA.n29 PRE_VLSA.n28 2.992
R4947 PRE_VLSA.n34 PRE_VLSA.n33 2.992
R4948 PRE_VLSA.n39 PRE_VLSA.n38 2.992
R4949 PRE_VLSA.n44 PRE_VLSA.n43 2.992
R4950 PRE_VLSA.n49 PRE_VLSA.n48 2.992
R4951 PRE_VLSA.n54 PRE_VLSA.n53 2.992
R4952 PRE_VLSA.n59 PRE_VLSA.n58 2.992
R4953 PRE_VLSA.n64 PRE_VLSA.n63 2.992
R4954 PRE_VLSA.n69 PRE_VLSA.n68 2.992
R4955 PRE_VLSA.n74 PRE_VLSA.n73 2.992
R4956 PRE_VLSA.n79 PRE_VLSA.n78 2.992
R4957 PRE_VLSA.n84 PRE_VLSA.n83 2.992
R4958 PRE_VLSA.n89 PRE_VLSA.n88 2.992
R4959 PRE_VLSA.n94 PRE_VLSA.n93 2.992
R4960 PRE_VLSA.n99 PRE_VLSA.n98 2.992
R4961 PRE_VLSA.n104 PRE_VLSA.n103 2.992
R4962 PRE_VLSA.n109 PRE_VLSA.n108 2.992
R4963 PRE_VLSA.n114 PRE_VLSA.n113 2.992
R4964 PRE_VLSA.n119 PRE_VLSA.n118 2.992
R4965 PRE_VLSA.n124 PRE_VLSA.n123 2.992
R4966 PRE_VLSA.n129 PRE_VLSA.n128 2.992
R4967 PRE_VLSA.n134 PRE_VLSA.n133 2.992
R4968 PRE_VLSA.n139 PRE_VLSA.n138 2.992
R4969 PRE_VLSA.n144 PRE_VLSA.n143 2.992
R4970 PRE_VLSA.n149 PRE_VLSA.n148 2.992
R4971 PRE_VLSA.n154 PRE_VLSA.n153 2.246
R4972 PRE_VLSA.n6 PRE_VLSA.n5 1.635
R4973 PRE_VLSA.n16 PRE_VLSA.n15 1.635
R4974 PRE_VLSA.n26 PRE_VLSA.n25 1.635
R4975 PRE_VLSA.n36 PRE_VLSA.n35 1.635
R4976 PRE_VLSA.n46 PRE_VLSA.n45 1.635
R4977 PRE_VLSA.n56 PRE_VLSA.n55 1.635
R4978 PRE_VLSA.n66 PRE_VLSA.n65 1.635
R4979 PRE_VLSA.n76 PRE_VLSA.n75 1.635
R4980 PRE_VLSA.n86 PRE_VLSA.n85 1.635
R4981 PRE_VLSA.n96 PRE_VLSA.n95 1.635
R4982 PRE_VLSA.n106 PRE_VLSA.n105 1.635
R4983 PRE_VLSA.n116 PRE_VLSA.n115 1.635
R4984 PRE_VLSA.n126 PRE_VLSA.n125 1.635
R4985 PRE_VLSA.n136 PRE_VLSA.n135 1.635
R4986 PRE_VLSA.n146 PRE_VLSA.n145 1.635
R4987 PRE_VLSA.n5 PRE_VLSA.n4 0.041
R4988 PRE_VLSA.n10 PRE_VLSA.n9 0.041
R4989 PRE_VLSA.n15 PRE_VLSA.n14 0.041
R4990 PRE_VLSA.n20 PRE_VLSA.n19 0.041
R4991 PRE_VLSA.n25 PRE_VLSA.n24 0.041
R4992 PRE_VLSA.n30 PRE_VLSA.n29 0.041
R4993 PRE_VLSA.n35 PRE_VLSA.n34 0.041
R4994 PRE_VLSA.n40 PRE_VLSA.n39 0.041
R4995 PRE_VLSA.n45 PRE_VLSA.n44 0.041
R4996 PRE_VLSA.n50 PRE_VLSA.n49 0.041
R4997 PRE_VLSA.n55 PRE_VLSA.n54 0.041
R4998 PRE_VLSA.n60 PRE_VLSA.n59 0.041
R4999 PRE_VLSA.n65 PRE_VLSA.n64 0.041
R5000 PRE_VLSA.n70 PRE_VLSA.n69 0.041
R5001 PRE_VLSA.n75 PRE_VLSA.n74 0.041
R5002 PRE_VLSA.n80 PRE_VLSA.n79 0.041
R5003 PRE_VLSA.n85 PRE_VLSA.n84 0.041
R5004 PRE_VLSA.n90 PRE_VLSA.n89 0.041
R5005 PRE_VLSA.n95 PRE_VLSA.n94 0.041
R5006 PRE_VLSA.n100 PRE_VLSA.n99 0.041
R5007 PRE_VLSA.n105 PRE_VLSA.n104 0.041
R5008 PRE_VLSA.n110 PRE_VLSA.n109 0.041
R5009 PRE_VLSA.n115 PRE_VLSA.n114 0.041
R5010 PRE_VLSA.n120 PRE_VLSA.n119 0.041
R5011 PRE_VLSA.n125 PRE_VLSA.n124 0.041
R5012 PRE_VLSA.n130 PRE_VLSA.n129 0.041
R5013 PRE_VLSA.n135 PRE_VLSA.n134 0.041
R5014 PRE_VLSA.n140 PRE_VLSA.n139 0.041
R5015 PRE_VLSA.n145 PRE_VLSA.n144 0.041
R5016 PRE_VLSA.n150 PRE_VLSA.n149 0.041
R5017 PRE_VLSA.n154 PRE_VLSA.n151 0.041
R5018 PRE_VLSA.n155 PRE_VLSA.n154 0.041
R5019 PRE_VLSA.n149 PRE_VLSA.n146 0.021
R5020 PRE_VLSA.n144 PRE_VLSA.n141 0.021
R5021 PRE_VLSA.n139 PRE_VLSA.n136 0.021
R5022 PRE_VLSA.n134 PRE_VLSA.n131 0.021
R5023 PRE_VLSA.n129 PRE_VLSA.n126 0.021
R5024 PRE_VLSA.n124 PRE_VLSA.n121 0.021
R5025 PRE_VLSA.n119 PRE_VLSA.n116 0.021
R5026 PRE_VLSA.n114 PRE_VLSA.n111 0.021
R5027 PRE_VLSA.n109 PRE_VLSA.n106 0.021
R5028 PRE_VLSA.n104 PRE_VLSA.n101 0.021
R5029 PRE_VLSA.n99 PRE_VLSA.n96 0.021
R5030 PRE_VLSA.n94 PRE_VLSA.n91 0.021
R5031 PRE_VLSA.n89 PRE_VLSA.n86 0.021
R5032 PRE_VLSA.n84 PRE_VLSA.n81 0.021
R5033 PRE_VLSA.n79 PRE_VLSA.n76 0.021
R5034 PRE_VLSA.n74 PRE_VLSA.n71 0.021
R5035 PRE_VLSA.n69 PRE_VLSA.n66 0.021
R5036 PRE_VLSA.n64 PRE_VLSA.n61 0.021
R5037 PRE_VLSA.n59 PRE_VLSA.n56 0.021
R5038 PRE_VLSA.n54 PRE_VLSA.n51 0.021
R5039 PRE_VLSA.n49 PRE_VLSA.n46 0.021
R5040 PRE_VLSA.n44 PRE_VLSA.n41 0.021
R5041 PRE_VLSA.n39 PRE_VLSA.n36 0.021
R5042 PRE_VLSA.n34 PRE_VLSA.n31 0.021
R5043 PRE_VLSA.n29 PRE_VLSA.n26 0.021
R5044 PRE_VLSA.n24 PRE_VLSA.n21 0.021
R5045 PRE_VLSA.n19 PRE_VLSA.n16 0.021
R5046 PRE_VLSA.n14 PRE_VLSA.n11 0.021
R5047 PRE_VLSA.n9 PRE_VLSA.n6 0.021
R5048 PRE_VLSA.n4 PRE_VLSA.n1 0.021
R5049 PRE_VLSA.n3 PRE_VLSA.n2 0.014
R5050 PRE_VLSA.n8 PRE_VLSA.n7 0.014
R5051 PRE_VLSA.n13 PRE_VLSA.n12 0.014
R5052 PRE_VLSA.n18 PRE_VLSA.n17 0.014
R5053 PRE_VLSA.n23 PRE_VLSA.n22 0.014
R5054 PRE_VLSA.n28 PRE_VLSA.n27 0.014
R5055 PRE_VLSA.n33 PRE_VLSA.n32 0.014
R5056 PRE_VLSA.n38 PRE_VLSA.n37 0.014
R5057 PRE_VLSA.n43 PRE_VLSA.n42 0.014
R5058 PRE_VLSA.n48 PRE_VLSA.n47 0.014
R5059 PRE_VLSA.n53 PRE_VLSA.n52 0.014
R5060 PRE_VLSA.n58 PRE_VLSA.n57 0.014
R5061 PRE_VLSA.n63 PRE_VLSA.n62 0.014
R5062 PRE_VLSA.n68 PRE_VLSA.n67 0.014
R5063 PRE_VLSA.n73 PRE_VLSA.n72 0.014
R5064 PRE_VLSA.n78 PRE_VLSA.n77 0.014
R5065 PRE_VLSA.n83 PRE_VLSA.n82 0.014
R5066 PRE_VLSA.n88 PRE_VLSA.n87 0.014
R5067 PRE_VLSA.n93 PRE_VLSA.n92 0.014
R5068 PRE_VLSA.n98 PRE_VLSA.n97 0.014
R5069 PRE_VLSA.n103 PRE_VLSA.n102 0.014
R5070 PRE_VLSA.n108 PRE_VLSA.n107 0.014
R5071 PRE_VLSA.n113 PRE_VLSA.n112 0.014
R5072 PRE_VLSA.n118 PRE_VLSA.n117 0.014
R5073 PRE_VLSA.n123 PRE_VLSA.n122 0.014
R5074 PRE_VLSA.n128 PRE_VLSA.n127 0.014
R5075 PRE_VLSA.n133 PRE_VLSA.n132 0.014
R5076 PRE_VLSA.n138 PRE_VLSA.n137 0.014
R5077 PRE_VLSA.n143 PRE_VLSA.n142 0.014
R5078 PRE_VLSA.n148 PRE_VLSA.n147 0.014
R5079 PRE_VLSA.n153 PRE_VLSA.n152 0.011
R5080 VDD.t555 VDD.t1221 1134.86
R5081 VDD.t1003 VDD.t2165 1028.47
R5082 VDD.t943 VDD.t491 970.652
R5083 VDD.t977 VDD.t2163 970.652
R5084 VDD.t28 VDD.t1604 970.652
R5085 VDD.t338 VDD.t1965 970.652
R5086 VDD.t879 VDD.t473 970.652
R5087 VDD.t1506 VDD.t535 970.652
R5088 VDD.t1883 VDD.t1747 970.652
R5089 VDD.t1022 VDD.t841 970.652
R5090 VDD.t2007 VDD.t1852 970.652
R5091 VDD.t461 VDD.t937 970.652
R5092 VDD.t2282 VDD.t453 970.652
R5093 VDD.t967 VDD.t547 970.652
R5094 VDD.t2204 VDD.t971 970.652
R5095 VDD.t1969 VDD.t793 970.652
R5096 VDD.t1700 VDD.t2262 970.652
R5097 VDD.t766 VDD.t2202 970.652
R5098 VDD.t384 VDD.t1243 970.652
R5099 VDD.t1877 VDD.t2005 970.652
R5100 VDD.t1939 VDD.t2145 970.652
R5101 VDD.t521 VDD.t1387 970.652
R5102 VDD.t1482 VDD.t1184 970.652
R5103 VDD.t883 VDD.t2179 970.652
R5104 VDD.t2175 VDD.t2237 970.652
R5105 VDD.t2224 VDD.t1799 970.652
R5106 VDD.t439 VDD.t780 970.652
R5107 VDD.t1170 VDD.t437 970.652
R5108 VDD.t1635 VDD.t553 970.652
R5109 VDD.t2141 VDD.t1941 970.652
R5110 VDD.t727 VDD.t58 970.652
R5111 VDD.t2157 VDD.t774 970.652
R5112 VDD.t1973 VDD.t2159 970.652
R5113 VDD.t1474 VDD.t1458 970.652
R5114 VDD.t1464 VDD.t993 970.652
R5115 VDD.t709 VDD.t2139 970.652
R5116 VDD.t503 VDD.t1702 970.652
R5117 VDD.t1311 VDD.t34 970.652
R5118 VDD.t609 VDD.t917 970.652
R5119 VDD.t1943 VDD.t433 970.652
R5120 VDD.t1048 VDD.t8 970.652
R5121 VDD.t20 VDD.t1561 970.652
R5122 VDD.t1631 VDD.t1706 970.652
R5123 VDD.t651 VDD.t1557 970.652
R5124 VDD.t1690 VDD.t1520 970.652
R5125 VDD.t711 VDD.t2131 970.652
R5126 VDD.t1016 VDD.t368 970.652
R5127 VDD.t44 VDD.t1080 970.652
R5128 VDD.t2274 VDD.t48 970.652
R5129 VDD.t1355 VDD.t829 970.652
R5130 VDD.t961 VDD.t667 970.652
R5131 VDD.t2246 VDD.t455 970.652
R5132 VDD.t981 VDD.t1818 970.652
R5133 VDD.t1247 VDD.t1842 970.652
R5134 VDD.t1696 VDD.t748 970.652
R5135 VDD.t1309 VDD.t1229 970.652
R5136 VDD.t669 VDD.t1719 970.652
R5137 VDD.t1911 VDD.t1812 970.652
R5138 VDD.t607 VDD.t380 970.652
R5139 VDD.t795 VDD.t1625 970.652
R5140 VDD.t1987 VDD.t807 970.652
R5141 VDD.t617 VDD.t2248 970.652
R5142 VDD.t2135 VDD.t891 970.652
R5143 VDD.t647 VDD.t1496 970.652
R5144 VDD.t1657 VDD.t649 970.652
R5145 VDD.t531 VDD.t1623 970.652
R5146 VDD.t1343 VDD.t1034 970.652
R5147 VDD.t579 VDD.t1369 970.652
R5148 VDD.t1584 VDD.t1397 970.652
R5149 VDD.t409 VDD.t1492 970.652
R5150 VDD.t931 VDD.t2101 970.652
R5151 VDD.t26 VDD.t1838 970.652
R5152 VDD.t758 VDD.t969 970.652
R5153 VDD.t1858 VDD.t1423 970.652
R5154 VDD.t1565 VDD.t392 970.652
R5155 VDD.t1327 VDD.t799 970.652
R5156 VDD.t459 VDD.t760 970.652
R5157 VDD.t2099 VDD.t1830 970.652
R5158 VDD.t786 VDD.t52 970.652
R5159 VDD.t725 VDD.t1735 970.652
R5160 VDD.t778 VDD.t770 970.652
R5161 VDD.t1721 VDD.t1759 970.652
R5162 VDD.t2200 VDD.t2107 970.652
R5163 VDD.t1686 VDD.t1494 970.652
R5164 VDD.t447 VDD.t390 970.652
R5165 VDD.t376 VDD.t939 970.652
R5166 VDD.t559 VDD.t1753 970.652
R5167 VDD.t481 VDD.t1266 970.652
R5168 VDD.t2169 VDD.t1715 970.652
R5169 VDD.t1713 VDD.t1543 970.652
R5170 VDD.t1959 VDD.t66 970.652
R5171 VDD.t12 VDD.t1953 970.652
R5172 VDD.t1761 VDD.t2171 970.652
R5173 VDD.t1361 VDD.t1297 970.652
R5174 VDD.t1299 VDD.t1359 970.652
R5175 VDD.t615 VDD.t911 970.652
R5176 VDD.t729 VDD.t2161 970.652
R5177 VDD.t70 VDD.t2184 970.652
R5178 VDD.t2206 VDD.t1606 970.652
R5179 VDD.t1572 VDD.t1188 970.652
R5180 VDD.t837 VDD.t1331 970.652
R5181 VDD.t1680 VDD.t1541 970.652
R5182 VDD.t991 VDD.t959 970.652
R5183 VDD.t853 VDD.t907 970.652
R5184 VDD.t1249 VDD.t465 970.652
R5185 VDD.t507 VDD.t1611 970.652
R5186 VDD.t1594 VDD.t2149 970.652
R5187 VDD.t2188 VDD.t589 970.652
R5188 VDD.t2121 VDD.t40 970.652
R5189 VDD.t2115 VDD.t1377 970.652
R5190 VDD.t951 VDD.t1028 970.652
R5191 VDD.t1313 VDD.t605 970.652
R5192 VDD.t661 VDD.t683 970.652
R5193 VDD.t1929 VDD.t2212 970.652
R5194 VDD.t673 VDD.t583 970.652
R5195 VDD.t689 VDD.t2220 970.652
R5196 VDD.t2210 VDD.t2186 970.652
R5197 VDD.t1767 VDD.t2264 970.652
R5198 VDD.t1771 VDD.t889 970.652
R5199 VDD.t953 VDD.t516 970.652
R5200 VDD.t561 VDD.t360 970.652
R5201 VDD.t621 VDD.t1391 970.652
R5202 VDD.t519 VDD.t1895 970.652
R5203 VDD.t1476 VDD.t1885 970.652
R5204 VDD.t6 VDD.t1472 970.652
R5205 VDD.t46 VDD.t1100 970.652
R5206 VDD.t1102 VDD.t791 970.652
R5207 VDD.t1425 VDD.t1961 970.652
R5208 VDD.t2167 VDD.t1014 970.652
R5209 VDD.t1985 VDD.t2198 970.652
R5210 VDD.t1480 VDD.t1844 970.652
R5211 VDD.t413 VDD.t2173 970.652
R5212 VDD.t2268 VDD.t328 970.652
R5213 VDD.t1574 VDD.t1286 970.652
R5214 VDD.t627 VDD.t354 970.652
R5215 VDD.t1470 VDD.t1613 970.652
R5216 VDD.t1602 VDD.t318 970.652
R5217 VDD.t50 VDD.t955 970.652
R5218 VDD.t1820 VDD.t1539 970.652
R5219 VDD.t423 VDD.t1795 970.652
R5220 VDD.t1367 VDD.t1708 970.652
R5221 VDD.t457 VDD.t1801 970.652
R5222 VDD.t1803 VDD.t585 970.652
R5223 VDD.t2222 VDD.t1733 970.652
R5224 VDD.t312 VDD.t995 970.652
R5225 VDD.t601 VDD.t1921 970.652
R5226 VDD.t593 VDD.t1516 970.652
R5227 VDD.t1264 VDD.t1661 970.652
R5228 VDD.t1663 VDD.t1967 970.652
R5229 VDD.t1777 VDD.t80 970.652
R5230 VDD.t1907 VDD.t1769 970.652
R5231 VDD.t1586 VDD.t549 970.652
R5232 VDD.t577 VDD.t1828 970.652
R5233 VDD.t1615 VDD.t1058 970.652
R5234 VDD.t370 VDD.t1860 970.652
R5235 VDD.t527 VDD.t1731 970.652
R5236 VDD.t1647 VDD.t653 970.652
R5237 VDD.t2252 VDD.t441 970.652
R5238 VDD.t1737 VDD.t1935 970.652
R5239 VDD.t813 VDD.t42 970.652
R5240 VDD.t2153 VDD.t825 970.652
R5241 VDD.t983 VDD.t1913 970.652
R5242 VDD.t1268 VDD.t1563 970.652
R5243 VDD.t310 VDD.t869 970.652
R5244 VDD.t1873 VDD.t1741 970.652
R5245 VDD.t1989 VDD.t989 970.652
R5246 VDD.t857 VDD.t2001 970.652
R5247 VDD.t340 VDD.t875 970.652
R5248 VDD.t1704 VDD.t1512 970.652
R5249 VDD.t913 VDD.t1793 970.652
R5250 VDD.t1417 VDD.t2233 970.652
R5251 VDD.t388 VDD.t599 970.652
R5252 VDD.t1526 VDD.t467 970.652
R5253 VDD.t1651 VDD.t1225 970.652
R5254 VDD.t475 VDD.t1779 970.652
R5255 VDD.t1893 VDD.t999 970.652
R5256 VDD.t1347 VDD.t1897 970.652
R5257 VDD.t947 VDD.t1010 970.652
R5258 VDD.t1272 VDD.t449 970.652
R5259 VDD.t1598 VDD.t1743 970.652
R5260 VDD.t1864 VDD.t1090 970.652
R5261 VDD.t1488 VDD.t1836 970.652
R5262 VDD.t545 VDD.t1745 970.652
R5263 VDD.t1408 VDD.t1421 970.652
R5264 VDD.t1848 VDD.t1383 970.652
R5265 VDD.t1385 VDD.t493 970.652
R5266 VDD.t833 VDD.t945 970.652
R5267 VDD.t1305 VDD.t831 970.652
R5268 VDD.t705 VDD.t1280 970.652
R5269 VDD.t358 VDD.t1284 970.652
R5270 VDD.t330 VDD.t923 970.652
R5271 VDD.t1524 VDD.t1098 970.652
R5272 VDD.t1518 VDD.t1846 970.652
R5273 VDD.t523 VDD.t1951 970.652
R5274 VDD.t16 VDD.t809 970.652
R5275 VDD.t1751 VDD.t514 970.652
R5276 VDD.t533 VDD.t1020 970.652
R5277 VDD.t1824 VDD.t597 970.652
R5278 VDD.t415 VDD.t587 970.652
R5279 VDD.t754 VDD.t2113 970.652
R5280 VDD.t2111 VDD.t1891 970.652
R5281 VDD.t657 VDD.t1412 970.652
R5282 VDD.t819 VDD.t1339 970.652
R5283 VDD.t1627 VDD.t1826 970.652
R5284 VDD.t1292 VDD.t1231 970.652
R5285 VDD.t2235 VDD.t2190 970.652
R5286 VDD.t2208 VDD.t1975 970.652
R5287 VDD.t1321 VDD.t1468 970.652
R5288 VDD.t975 VDD.t1323 970.652
R5289 VDD.t1633 VDD.t1723 970.652
R5290 VDD.t469 VDD.t1502 970.652
R5291 VDD.t851 VDD.t342 970.652
R5292 VDD.t1092 VDD.t1414 970.652
R5293 VDD.t78 VDD.t1046 970.652
R5294 VDD.t1881 VDD.t332 970.652
R5295 VDD.t1694 VDD.t489 970.652
R5296 VDD.t887 VDD.t715 970.652
R5297 VDD.t717 VDD.t1729 970.652
R5298 VDD.t1062 VDD.t659 970.652
R5299 VDD.t1995 VDD.t731 970.652
R5300 VDD.t1931 VDD.t1871 970.652
R5301 VDD.t537 VDD.t1582 970.652
R5302 VDD.t573 VDD.t895 970.652
R5303 VDD.t645 VDD.t74 970.652
R5304 VDD.t613 VDD.t935 970.652
R5305 VDD.t1174 VDD.t1692 970.652
R5306 VDD.t1927 VDD.t1274 970.652
R5307 VDD.t957 VDD.t2133 970.652
R5308 VDD.t1991 VDD.t1949 970.652
R5309 VDD.t1437 VDD.t1899 970.652
R5310 VDD.t762 VDD.t643 970.652
R5311 VDD.t352 VDD.t1404 970.652
R5312 VDD.t679 VDD.t405 970.652
R5313 VDD.t417 VDD.t403 970.652
R5314 VDD.t1439 VDD.t1875 970.652
R5315 VDD.t324 VDD.t563 970.652
R5316 VDD.t1333 VDD.t322 970.652
R5317 VDD.t1993 VDD.t1528 970.652
R5318 VDD.t386 VDD.t1453 970.652
R5319 VDD.t2009 VDD.t677 970.652
R5320 VDD.t2137 VDD.t2280 970.652
R5321 VDD.t695 VDD.t823 970.652
R5322 VDD.t855 VDD.t2284 970.652
R5323 VDD.t1032 VDD.t1629 970.652
R5324 VDD.t927 VDD.t1365 970.652
R5325 VDD.t835 VDD.t1064 970.652
R5326 VDD.t1038 VDD.t863 970.652
R5327 VDD.t1917 VDD.t501 970.652
R5328 VDD.t1050 VDD.t1822 970.652
R5329 VDD.t1617 VDD.t479 970.652
R5330 VDD.t2127 VDD.t346 970.652
R5331 VDD.t1808 VDD.t1909 970.652
R5332 VDD.t901 VDD.t477 970.652
R5333 VDD.t739 VDD.t374 970.652
R5334 VDD.t372 VDD.t1094 970.652
R5335 VDD.t713 VDD.t2231 970.652
R5336 VDD.t1484 VDD.t1773 970.652
R5337 VDD.t2123 VDD.t2155 970.652
R5338 VDD.n1621 VDD.t2286 696.666
R5339 VDD.n1469 VDD.t1052 696.666
R5340 VDD.n1325 VDD.t859 696.666
R5341 VDD.n1181 VDD.t1765 696.666
R5342 VDD.n1037 VDD.t1856 696.666
R5343 VDD.n893 VDD.t625 696.666
R5344 VDD.n749 VDD.t1241 696.666
R5345 VDD.n601 VDD.t1003 696.666
R5346 VDD.n671 VDD.t1486 695.289
R5347 VDD.n743 VDD.t1905 695.289
R5348 VDD.n815 VDD.t2272 695.289
R5349 VDD.n887 VDD.t1669 695.289
R5350 VDD.n959 VDD.t1887 695.289
R5351 VDD.n1031 VDD.t1739 695.289
R5352 VDD.n1103 VDD.t1345 695.289
R5353 VDD.n1175 VDD.t2181 695.289
R5354 VDD.n1247 VDD.t314 695.289
R5355 VDD.n1319 VDD.t1933 695.289
R5356 VDD.n1391 VDD.t1755 695.289
R5357 VDD.n1463 VDD.t2 695.289
R5358 VDD.n1535 VDD.t1401 695.289
R5359 VDD.n614 VDD.t1901 695.289
R5360 VDD.n1615 VDD.t1999 695.289
R5361 VDD.n532 VDD.t1431 695.289
R5362 VDD.t491 VDD.t1410 688.405
R5363 VDD.t1086 VDD.t943 688.405
R5364 VDD.n733 VDD.t1086 688.405
R5365 VDD.t897 VDD.t977 688.405
R5366 VDD.t2163 VDD.t28 688.405
R5367 VDD.t1604 VDD.t1592 688.405
R5368 VDD.t1965 VDD.t2125 688.405
R5369 VDD.t473 VDD.t338 688.405
R5370 VDD.t1608 VDD.t879 688.405
R5371 VDD.n718 VDD.t1608 688.405
R5372 VDD.t1547 VDD.t1506 688.405
R5373 VDD.t535 VDD.t1883 688.405
R5374 VDD.t1747 VDD.t1022 688.405
R5375 VDD.t841 VDD.t1643 688.405
R5376 VDD.t1852 VDD.t768 688.405
R5377 VDD.t937 VDD.t2007 688.405
R5378 VDD.t453 VDD.t461 688.405
R5379 VDD.t2254 VDD.t2282 688.405
R5380 VDD.n700 VDD.t2254 688.405
R5381 VDD.t985 VDD.t967 688.405
R5382 VDD.t547 VDD.t2204 688.405
R5383 VDD.t971 VDD.t973 688.405
R5384 VDD.t2262 VDD.t1969 688.405
R5385 VDD.t1486 VDD.t1700 688.405
R5386 VDD.t1840 VDD.t766 688.405
R5387 VDD.t2202 VDD.t784 688.405
R5388 VDD.t1243 VDD.t569 688.405
R5389 VDD.t1621 VDD.t384 688.405
R5390 VDD.n805 VDD.t1621 688.405
R5391 VDD.t1879 VDD.t1877 688.405
R5392 VDD.t2005 VDD.t1939 688.405
R5393 VDD.t2145 VDD.t2151 688.405
R5394 VDD.t1387 VDD.t411 688.405
R5395 VDD.t1184 VDD.t521 688.405
R5396 VDD.t764 VDD.t1482 688.405
R5397 VDD.n790 VDD.t764 688.405
R5398 VDD.t350 VDD.t883 688.405
R5399 VDD.t2179 VDD.t2175 688.405
R5400 VDD.t2237 VDD.t2224 688.405
R5401 VDD.t1799 VDD.t1168 688.405
R5402 VDD.t780 VDD.t776 688.405
R5403 VDD.t437 VDD.t439 688.405
R5404 VDD.t553 VDD.t1170 688.405
R5405 VDD.t1791 VDD.t1635 688.405
R5406 VDD.n772 VDD.t1791 688.405
R5407 VDD.t1427 VDD.t2141 688.405
R5408 VDD.t1941 VDD.t727 688.405
R5409 VDD.t58 VDD.t62 688.405
R5410 VDD.t2159 VDD.t2157 688.405
R5411 VDD.t1905 VDD.t1973 688.405
R5412 VDD.t1478 VDD.t1474 688.405
R5413 VDD.t1458 VDD.t1678 688.405
R5414 VDD.t993 VDD.t865 688.405
R5415 VDD.t721 VDD.t1464 688.405
R5416 VDD.n877 VDD.t721 688.405
R5417 VDD.t1903 VDD.t709 688.405
R5418 VDD.t2139 VDD.t503 688.405
R5419 VDD.t1702 VDD.t1257 688.405
R5420 VDD.t34 VDD.t24 688.405
R5421 VDD.t917 VDD.t1311 688.405
R5422 VDD.t1190 VDD.t609 688.405
R5423 VDD.n862 VDD.t1190 688.405
R5424 VDD.t2119 VDD.t1943 688.405
R5425 VDD.t433 VDD.t1048 688.405
R5426 VDD.t8 VDD.t20 688.405
R5427 VDD.t1561 VDD.t1012 688.405
R5428 VDD.t1706 VDD.t693 688.405
R5429 VDD.t1557 VDD.t1631 688.405
R5430 VDD.t1520 VDD.t651 688.405
R5431 VDD.t0 VDD.t1690 688.405
R5432 VDD.n844 VDD.t0 688.405
R5433 VDD.t701 VDD.t711 688.405
R5434 VDD.t2131 VDD.t1016 688.405
R5435 VDD.t368 VDD.t1007 688.405
R5436 VDD.t48 VDD.t44 688.405
R5437 VDD.t2272 VDD.t2274 688.405
R5438 VDD.t1357 VDD.t1355 688.405
R5439 VDD.t829 VDD.t1684 688.405
R5440 VDD.t667 VDD.t1866 688.405
R5441 VDD.t963 VDD.t961 688.405
R5442 VDD.n949 VDD.t963 688.405
R5443 VDD.t2226 VDD.t2246 688.405
R5444 VDD.t455 VDD.t981 688.405
R5445 VDD.t1818 VDD.t1329 688.405
R5446 VDD.t1842 VDD.t772 688.405
R5447 VDD.t748 VDD.t1247 688.405
R5448 VDD.t483 VDD.t1696 688.405
R5449 VDD.n934 VDD.t483 688.405
R5450 VDD.t1490 VDD.t1309 688.405
R5451 VDD.t1229 VDD.t669 688.405
R5452 VDD.t1719 VDD.t1911 688.405
R5453 VDD.t1812 VDD.t1282 688.405
R5454 VDD.t380 VDD.t529 688.405
R5455 VDD.t1625 VDD.t607 688.405
R5456 VDD.t807 VDD.t795 688.405
R5457 VDD.t2003 VDD.t1987 688.405
R5458 VDD.n916 VDD.t2003 688.405
R5459 VDD.t639 VDD.t617 688.405
R5460 VDD.t2248 VDD.t2135 688.405
R5461 VDD.t891 VDD.t782 688.405
R5462 VDD.t649 VDD.t647 688.405
R5463 VDD.t1669 VDD.t1657 688.405
R5464 VDD.t1325 VDD.t531 688.405
R5465 VDD.t1623 VDD.t1637 688.405
R5466 VDD.t1034 VDD.t344 688.405
R5467 VDD.t541 VDD.t1343 688.405
R5468 VDD.n1021 VDD.t541 688.405
R5469 VDD.t581 VDD.t579 688.405
R5470 VDD.t1369 VDD.t1584 688.405
R5471 VDD.t1397 VDD.t965 688.405
R5472 VDD.t1492 VDD.t671 688.405
R5473 VDD.t2101 VDD.t409 688.405
R5474 VDD.t2117 VDD.t931 688.405
R5475 VDD.n1006 VDD.t2117 688.405
R5476 VDD.t744 VDD.t26 688.405
R5477 VDD.t1838 VDD.t758 688.405
R5478 VDD.t969 VDD.t1858 688.405
R5479 VDD.t1423 VDD.t805 688.405
R5480 VDD.t392 VDD.t429 688.405
R5481 VDD.t799 VDD.t1565 688.405
R5482 VDD.t760 VDD.t1327 688.405
R5483 VDD.t1076 VDD.t459 688.405
R5484 VDD.n988 VDD.t1076 688.405
R5485 VDD.t2250 VDD.t2099 688.405
R5486 VDD.t1830 VDD.t786 688.405
R5487 VDD.t52 VDD.t38 688.405
R5488 VDD.t770 VDD.t725 688.405
R5489 VDD.t1887 VDD.t778 688.405
R5490 VDD.t1375 VDD.t1721 688.405
R5491 VDD.t1759 VDD.t443 688.405
R5492 VDD.t2107 VDD.t2256 688.405
R5493 VDD.t56 VDD.t2200 688.405
R5494 VDD.n1093 VDD.t56 688.405
R5495 VDD.t1717 VDD.t1686 688.405
R5496 VDD.t1494 VDD.t447 688.405
R5497 VDD.t390 VDD.t407 688.405
R5498 VDD.t939 VDD.t941 688.405
R5499 VDD.t1753 VDD.t376 688.405
R5500 VDD.t575 VDD.t559 688.405
R5501 VDD.n1078 VDD.t575 688.405
R5502 VDD.t451 VDD.t481 688.405
R5503 VDD.t1266 VDD.t2169 688.405
R5504 VDD.t1715 VDD.t1713 688.405
R5505 VDD.t1543 VDD.t14 688.405
R5506 VDD.t66 VDD.t82 688.405
R5507 VDD.t1953 VDD.t1959 688.405
R5508 VDD.t2171 VDD.t12 688.405
R5509 VDD.t1810 VDD.t1761 688.405
R5510 VDD.n1060 VDD.t1810 688.405
R5511 VDD.t1363 VDD.t1361 688.405
R5512 VDD.t1297 VDD.t1299 688.405
R5513 VDD.t1359 VDD.t435 688.405
R5514 VDD.t2161 VDD.t615 688.405
R5515 VDD.t1739 VDD.t729 688.405
R5516 VDD.t36 VDD.t70 688.405
R5517 VDD.t2184 VDD.t2177 688.405
R5518 VDD.t1606 VDD.t987 688.405
R5519 VDD.t2196 VDD.t2206 688.405
R5520 VDD.n1165 VDD.t2196 688.405
R5521 VDD.t1869 VDD.t1572 688.405
R5522 VDD.t1188 VDD.t837 688.405
R5523 VDD.t1331 VDD.t1278 688.405
R5524 VDD.t1541 VDD.t1259 688.405
R5525 VDD.t959 VDD.t1680 688.405
R5526 VDD.t867 VDD.t991 688.405
R5527 VDD.n1150 VDD.t867 688.405
R5528 VDD.t1785 VDD.t853 688.405
R5529 VDD.t907 VDD.t1249 688.405
R5530 VDD.t465 VDD.t507 688.405
R5531 VDD.t1611 VDD.t485 688.405
R5532 VDD.t2149 VDD.t320 688.405
R5533 VDD.t589 VDD.t1594 688.405
R5534 VDD.t40 VDD.t2188 688.405
R5535 VDD.t1862 VDD.t2121 688.405
R5536 VDD.n1132 VDD.t1862 688.405
R5537 VDD.t2103 VDD.t2115 688.405
R5538 VDD.t1377 VDD.t951 688.405
R5539 VDD.t1028 VDD.t1533 688.405
R5540 VDD.t683 VDD.t1313 688.405
R5541 VDD.t1345 VDD.t661 688.405
R5542 VDD.t54 VDD.t1929 688.405
R5543 VDD.t2212 VDD.t2218 688.405
R5544 VDD.t583 VDD.t1026 688.405
R5545 VDD.t675 VDD.t673 688.405
R5546 VDD.n1237 VDD.t675 688.405
R5547 VDD.t685 VDD.t689 688.405
R5548 VDD.t2220 VDD.t2210 688.405
R5549 VDD.t2186 VDD.t815 688.405
R5550 VDD.t2264 VDD.t2266 688.405
R5551 VDD.t889 VDD.t1767 688.405
R5552 VDD.t1373 VDD.t1771 688.405
R5553 VDD.n1222 VDD.t1373 688.405
R5554 VDD.t687 VDD.t953 688.405
R5555 VDD.t516 VDD.t561 688.405
R5556 VDD.t360 VDD.t621 688.405
R5557 VDD.t1391 VDD.t1303 688.405
R5558 VDD.t1895 VDD.t949 688.405
R5559 VDD.t1885 VDD.t519 688.405
R5560 VDD.t1472 VDD.t1476 688.405
R5561 VDD.t10 VDD.t6 688.405
R5562 VDD.n1204 VDD.t10 688.405
R5563 VDD.t84 VDD.t46 688.405
R5564 VDD.t1100 VDD.t1102 688.405
R5565 VDD.t791 VDD.t817 688.405
R5566 VDD.t1014 VDD.t1425 688.405
R5567 VDD.t2181 VDD.t2167 688.405
R5568 VDD.t1919 VDD.t1985 688.405
R5569 VDD.t2198 VDD.t2214 688.405
R5570 VDD.t1844 VDD.t463 688.405
R5571 VDD.t1816 VDD.t1480 688.405
R5572 VDD.n1309 VDD.t1816 688.405
R5573 VDD.t505 VDD.t413 688.405
R5574 VDD.t2173 VDD.t2268 688.405
R5575 VDD.t328 VDD.t2147 688.405
R5576 VDD.t1286 VDD.t2216 688.405
R5577 VDD.t354 VDD.t1574 688.405
R5578 VDD.t1569 VDD.t627 688.405
R5579 VDD.n1294 VDD.t1569 688.405
R5580 VDD.t1056 VDD.t1470 688.405
R5581 VDD.t1613 VDD.t1602 688.405
R5582 VDD.t318 VDD.t50 688.405
R5583 VDD.t955 VDD.t382 688.405
R5584 VDD.t1539 VDD.t595 688.405
R5585 VDD.t1795 VDD.t1820 688.405
R5586 VDD.t1708 VDD.t423 688.405
R5587 VDD.t925 VDD.t1367 688.405
R5588 VDD.n1276 VDD.t925 688.405
R5589 VDD.t1351 VDD.t457 688.405
R5590 VDD.t1801 VDD.t1803 688.405
R5591 VDD.t585 VDD.t655 688.405
R5592 VDD.t995 VDD.t2222 688.405
R5593 VDD.t314 VDD.t312 688.405
R5594 VDD.t603 VDD.t601 688.405
R5595 VDD.t1921 VDD.t1925 688.405
R5596 VDD.t1516 VDD.t1522 688.405
R5597 VDD.t1435 VDD.t593 688.405
R5598 VDD.n1381 VDD.t1435 688.405
R5599 VDD.t691 VDD.t1264 688.405
R5600 VDD.t1661 VDD.t1663 688.405
R5601 VDD.t1967 VDD.t2093 688.405
R5602 VDD.t80 VDD.t1659 688.405
R5603 VDD.t1769 VDD.t1777 688.405
R5604 VDD.t1971 VDD.t1907 688.405
R5605 VDD.n1366 VDD.t1971 688.405
R5606 VDD.t567 VDD.t1586 688.405
R5607 VDD.t549 VDD.t577 688.405
R5608 VDD.t1828 VDD.t1615 688.405
R5609 VDD.t1058 VDD.t1588 688.405
R5610 VDD.t1860 VDD.t641 688.405
R5611 VDD.t1731 VDD.t370 688.405
R5612 VDD.t653 VDD.t527 688.405
R5613 VDD.t1649 VDD.t1647 688.405
R5614 VDD.n1348 VDD.t1649 688.405
R5615 VDD.t756 VDD.t2252 688.405
R5616 VDD.t441 VDD.t1737 688.405
R5617 VDD.t1935 VDD.t1937 688.405
R5618 VDD.t825 VDD.t813 688.405
R5619 VDD.t1933 VDD.t2153 688.405
R5620 VDD.t1395 VDD.t983 688.405
R5621 VDD.t1913 VDD.t2143 688.405
R5622 VDD.t1563 VDD.t495 688.405
R5623 VDD.t707 VDD.t1268 688.405
R5624 VDD.n1453 VDD.t707 688.405
R5625 VDD.t316 VDD.t310 688.405
R5626 VDD.t869 VDD.t1873 688.405
R5627 VDD.t1741 VDD.t1545 688.405
R5628 VDD.t989 VDD.t487 688.405
R5629 VDD.t2001 VDD.t1989 688.405
R5630 VDD.t1783 VDD.t857 688.405
R5631 VDD.n1438 VDD.t1783 688.405
R5632 VDD.t1261 VDD.t340 688.405
R5633 VDD.t875 VDD.t1704 688.405
R5634 VDD.t1512 VDD.t913 688.405
R5635 VDD.t1793 VDD.t1460 688.405
R5636 VDD.t2233 VDD.t2241 688.405
R5637 VDD.t599 VDD.t1417 688.405
R5638 VDD.t467 VDD.t388 688.405
R5639 VDD.t525 VDD.t1526 688.405
R5640 VDD.n1420 VDD.t525 688.405
R5641 VDD.t591 VDD.t1651 688.405
R5642 VDD.t1225 VDD.t475 688.405
R5643 VDD.t1779 VDD.t885 688.405
R5644 VDD.t1897 VDD.t1893 688.405
R5645 VDD.t1755 VDD.t1347 688.405
R5646 VDD.t399 VDD.t947 688.405
R5647 VDD.t1010 VDD.t539 688.405
R5648 VDD.t449 VDD.t1379 688.405
R5649 VDD.t750 VDD.t1272 688.405
R5650 VDD.n1525 VDD.t750 688.405
R5651 VDD.t1042 VDD.t1598 688.405
R5652 VDD.t1743 VDD.t1864 688.405
R5653 VDD.t1090 VDD.t903 688.405
R5654 VDD.t1836 VDD.t1688 688.405
R5655 VDD.t1745 VDD.t1488 688.405
R5656 VDD.t1233 VDD.t545 688.405
R5657 VDD.n1510 VDD.t1233 688.405
R5658 VDD.t1406 VDD.t1408 688.405
R5659 VDD.t1421 VDD.t1848 688.405
R5660 VDD.t1383 VDD.t1385 688.405
R5661 VDD.t493 VDD.t1559 688.405
R5662 VDD.t945 VDD.t1578 688.405
R5663 VDD.t831 VDD.t833 688.405
R5664 VDD.t1280 VDD.t1305 688.405
R5665 VDD.t611 VDD.t705 688.405
R5666 VDD.n1492 VDD.t611 688.405
R5667 VDD.t933 VDD.t358 688.405
R5668 VDD.t1284 VDD.t330 688.405
R5669 VDD.t923 VDD.t1665 688.405
R5670 VDD.t1846 VDD.t1524 688.405
R5671 VDD.t2 VDD.t1518 688.405
R5672 VDD.t1178 VDD.t523 688.405
R5673 VDD.t1951 VDD.t2129 688.405
R5674 VDD.t809 VDD.t735 688.405
R5675 VDD.t2192 VDD.t16 688.405
R5676 VDD.n1597 VDD.t2192 688.405
R5677 VDD.t1186 VDD.t1751 688.405
R5678 VDD.t514 VDD.t533 688.405
R5679 VDD.t1020 VDD.t1024 688.405
R5680 VDD.t597 VDD.t1555 688.405
R5681 VDD.t587 VDD.t1824 688.405
R5682 VDD.t921 VDD.t415 688.405
R5683 VDD.n1582 VDD.t921 688.405
R5684 VDD.t1498 VDD.t754 688.405
R5685 VDD.t2113 VDD.t2111 688.405
R5686 VDD.t1891 VDD.t657 688.405
R5687 VDD.t1412 VDD.t378 688.405
R5688 VDD.t1339 VDD.t1341 688.405
R5689 VDD.t1826 VDD.t819 688.405
R5690 VDD.t1231 VDD.t1627 688.405
R5691 VDD.t499 VDD.t1292 688.405
R5692 VDD.n1564 VDD.t499 688.405
R5693 VDD.t881 VDD.t2235 688.405
R5694 VDD.t2190 VDD.t2208 688.405
R5695 VDD.t1975 VDD.t929 688.405
R5696 VDD.t1323 VDD.t1321 688.405
R5697 VDD.t1401 VDD.t975 688.405
R5698 VDD.t1500 VDD.t1633 688.405
R5699 VDD.t1723 VDD.t1725 688.405
R5700 VDD.t1502 VDD.t801 688.405
R5701 VDD.t1641 VDD.t469 688.405
R5702 VDD.n661 VDD.t1641 688.405
R5703 VDD.t1667 VDD.t851 688.405
R5704 VDD.t342 VDD.t1092 688.405
R5705 VDD.t1414 VDD.t909 688.405
R5706 VDD.t1046 VDD.t629 688.405
R5707 VDD.t332 VDD.t78 688.405
R5708 VDD.t1854 VDD.t1881 688.405
R5709 VDD.n646 VDD.t1854 688.405
R5710 VDD.t905 VDD.t1694 688.405
R5711 VDD.t489 VDD.t887 688.405
R5712 VDD.t715 VDD.t717 688.405
R5713 VDD.t1729 VDD.t1963 688.405
R5714 VDD.t659 VDD.t1915 688.405
R5715 VDD.t731 VDD.t1062 688.405
R5716 VDD.t1871 VDD.t1995 688.405
R5717 VDD.t1923 VDD.t1931 688.405
R5718 VDD.n628 VDD.t1923 688.405
R5719 VDD.t1040 VDD.t537 688.405
R5720 VDD.t1582 VDD.t573 688.405
R5721 VDD.t895 VDD.t1682 688.405
R5722 VDD.t935 VDD.t645 688.405
R5723 VDD.t1901 VDD.t613 688.405
R5724 VDD.t1957 VDD.t1174 688.405
R5725 VDD.t1692 VDD.t697 688.405
R5726 VDD.t1274 VDD.t631 688.405
R5727 VDD.t1983 VDD.t1927 688.405
R5728 VDD.n1608 VDD.t1983 688.405
R5729 VDD.t1576 VDD.t957 688.405
R5730 VDD.t2133 VDD.t1991 688.405
R5731 VDD.t1949 VDD.t1945 688.405
R5732 VDD.t1899 VDD.t2097 688.405
R5733 VDD.t643 VDD.t1437 688.405
R5734 VDD.t445 VDD.t762 688.405
R5735 VDD.n1610 VDD.t445 688.405
R5736 VDD.t1074 VDD.t352 688.405
R5737 VDD.t1404 VDD.t679 688.405
R5738 VDD.t405 VDD.t417 688.405
R5739 VDD.t403 VDD.t395 688.405
R5740 VDD.t1875 VDD.t1239 688.405
R5741 VDD.t563 VDD.t1439 688.405
R5742 VDD.t322 VDD.t324 688.405
R5743 VDD.t843 VDD.t1333 688.405
R5744 VDD.n1612 VDD.t843 688.405
R5745 VDD.t2243 VDD.t1993 688.405
R5746 VDD.t1528 VDD.t386 688.405
R5747 VDD.t1453 VDD.t1671 688.405
R5748 VDD.t2280 VDD.t2009 688.405
R5749 VDD.t1999 VDD.t2137 688.405
R5750 VDD.t557 VDD.t695 688.405
R5751 VDD.t823 VDD.t821 688.405
R5752 VDD.t2284 VDD.t1393 688.405
R5753 VDD.t1066 VDD.t855 688.405
R5754 VDD.n589 VDD.t1066 688.405
R5755 VDD.t1781 VDD.t1032 688.405
R5756 VDD.t1629 VDD.t927 688.405
R5757 VDD.t1365 VDD.t839 688.405
R5758 VDD.t1064 VDD.t703 688.405
R5759 VDD.t863 VDD.t835 688.405
R5760 VDD.t1301 VDD.t1038 688.405
R5761 VDD.n527 VDD.t1301 688.405
R5762 VDD.t1551 VDD.t1917 688.405
R5763 VDD.t501 VDD.t1050 688.405
R5764 VDD.t1822 VDD.t1617 688.405
R5765 VDD.t479 VDD.t356 688.405
R5766 VDD.t346 VDD.t1889 688.405
R5767 VDD.t1909 VDD.t2127 688.405
R5768 VDD.t477 VDD.t1808 688.405
R5769 VDD.t421 VDD.t901 688.405
R5770 VDD.n529 VDD.t421 688.405
R5771 VDD.t737 VDD.t739 688.405
R5772 VDD.t374 VDD.t372 688.405
R5773 VDD.t1094 VDD.t1389 688.405
R5774 VDD.t1773 VDD.t713 688.405
R5775 VDD.t1431 VDD.t1484 688.405
R5776 VDD.t1947 VDD.t2123 688.405
R5777 VDD.t2155 VDD.t2228 688.405
R5778 VDD.t793 VDD.t1757 681.521
R5779 VDD.n671 VDD.t1840 681.521
R5780 VDD.t774 VDD.t633 681.521
R5781 VDD.n743 VDD.t1478 681.521
R5782 VDD.t1080 VDD.t1078 681.521
R5783 VDD.n815 VDD.t1357 681.521
R5784 VDD.t1496 VDD.t1462 681.521
R5785 VDD.n887 VDD.t1325 681.521
R5786 VDD.t1735 VDD.t1514 681.521
R5787 VDD.n959 VDD.t1375 681.521
R5788 VDD.t911 VDD.t1245 681.521
R5789 VDD.n1031 VDD.t36 681.521
R5790 VDD.t605 VDD.t1255 681.521
R5791 VDD.n1103 VDD.t54 681.521
R5792 VDD.t1961 VDD.t1955 681.521
R5793 VDD.n1175 VDD.t1919 681.521
R5794 VDD.t1733 VDD.t1805 681.521
R5795 VDD.n1247 VDD.t603 681.521
R5796 VDD.t42 VDD.t64 681.521
R5797 VDD.n1319 VDD.t1395 681.521
R5798 VDD.t999 VDD.t1001 681.521
R5799 VDD.n1391 VDD.t399 681.521
R5800 VDD.t1098 VDD.t733 681.521
R5801 VDD.n1463 VDD.t1178 681.521
R5802 VDD.t1468 VDD.t1349 681.521
R5803 VDD.n1535 VDD.t1500 681.521
R5804 VDD.t74 VDD.t68 681.521
R5805 VDD.n614 VDD.t1957 681.521
R5806 VDD.t677 VDD.t899 681.521
R5807 VDD.n1615 VDD.t557 681.521
R5808 VDD.t2231 VDD.t2239 681.521
R5809 VDD.n532 VDD.t1947 681.521
R5810 VDD.n733 VDD.t897 667.753
R5811 VDD.n805 VDD.t1879 667.753
R5812 VDD.n877 VDD.t1903 667.753
R5813 VDD.n949 VDD.t2226 667.753
R5814 VDD.n1021 VDD.t581 667.753
R5815 VDD.n1093 VDD.t1717 667.753
R5816 VDD.n1165 VDD.t1869 667.753
R5817 VDD.n1237 VDD.t685 667.753
R5818 VDD.n1309 VDD.t505 667.753
R5819 VDD.n1381 VDD.t691 667.753
R5820 VDD.n1453 VDD.t316 667.753
R5821 VDD.n1525 VDD.t1042 667.753
R5822 VDD.n1597 VDD.t1186 667.753
R5823 VDD.n661 VDD.t1667 667.753
R5824 VDD.n1608 VDD.t1576 667.753
R5825 VDD.n589 VDD.t1781 667.753
R5826 VDD.n1621 VDD.t555 633.333
R5827 VDD.n1469 VDD.t2091 633.333
R5828 VDD.n1325 VDD.t803 633.333
R5829 VDD.n1181 VDD.t497 633.333
R5830 VDD.n1037 VDD.t873 633.333
R5831 VDD.n893 VDD.t510 633.333
R5832 VDD.n749 VDD.t1251 633.333
R5833 VDD.n601 VDD.t637 633.333
R5834 VDD.t1410 VDD.n732 612.681
R5835 VDD.t569 VDD.n804 612.681
R5836 VDD.t865 VDD.n876 612.681
R5837 VDD.t1866 VDD.n948 612.681
R5838 VDD.t344 VDD.n1020 612.681
R5839 VDD.t2256 VDD.n1092 612.681
R5840 VDD.t987 VDD.n1164 612.681
R5841 VDD.t1026 VDD.n1236 612.681
R5842 VDD.t463 VDD.n1308 612.681
R5843 VDD.t1522 VDD.n1380 612.681
R5844 VDD.t495 VDD.n1452 612.681
R5845 VDD.t1379 VDD.n1524 612.681
R5846 VDD.t735 VDD.n1596 612.681
R5847 VDD.t801 VDD.n660 612.681
R5848 VDD.t631 VDD.n1607 612.681
R5849 VDD.t1393 VDD.n588 612.681
R5850 VDD.n700 VDD.t985 564.492
R5851 VDD.t784 VDD.n670 564.492
R5852 VDD.n772 VDD.t1427 564.492
R5853 VDD.t1678 VDD.n742 564.492
R5854 VDD.n844 VDD.t701 564.492
R5855 VDD.t1684 VDD.n814 564.492
R5856 VDD.n916 VDD.t639 564.492
R5857 VDD.t1637 VDD.n886 564.492
R5858 VDD.n988 VDD.t2250 564.492
R5859 VDD.t443 VDD.n958 564.492
R5860 VDD.n1060 VDD.t1363 564.492
R5861 VDD.t2177 VDD.n1030 564.492
R5862 VDD.n1132 VDD.t2103 564.492
R5863 VDD.t2218 VDD.n1102 564.492
R5864 VDD.n1204 VDD.t84 564.492
R5865 VDD.t2214 VDD.n1174 564.492
R5866 VDD.n1276 VDD.t1351 564.492
R5867 VDD.t1925 VDD.n1246 564.492
R5868 VDD.n1348 VDD.t756 564.492
R5869 VDD.t2143 VDD.n1318 564.492
R5870 VDD.n1420 VDD.t591 564.492
R5871 VDD.t539 VDD.n1390 564.492
R5872 VDD.n1492 VDD.t933 564.492
R5873 VDD.t2129 VDD.n1462 564.492
R5874 VDD.n1564 VDD.t881 564.492
R5875 VDD.t1725 VDD.n1534 564.492
R5876 VDD.n628 VDD.t1040 564.492
R5877 VDD.t697 VDD.n613 564.492
R5878 VDD.n1612 VDD.t2243 564.492
R5879 VDD.t821 VDD.n1614 564.492
R5880 VDD.n529 VDD.t737 564.492
R5881 VDD.t2228 VDD.n531 564.492
R5882 VDD.n718 VDD.t1547 557.608
R5883 VDD.n790 VDD.t350 557.608
R5884 VDD.n862 VDD.t2119 557.608
R5885 VDD.n934 VDD.t1490 557.608
R5886 VDD.n1006 VDD.t744 557.608
R5887 VDD.n1078 VDD.t451 557.608
R5888 VDD.n1150 VDD.t1785 557.608
R5889 VDD.n1222 VDD.t687 557.608
R5890 VDD.n1294 VDD.t1056 557.608
R5891 VDD.n1366 VDD.t567 557.608
R5892 VDD.n1438 VDD.t1261 557.608
R5893 VDD.n1510 VDD.t1406 557.608
R5894 VDD.n1582 VDD.t1498 557.608
R5895 VDD.n646 VDD.t905 557.608
R5896 VDD.n1610 VDD.t1074 557.608
R5897 VDD.n527 VDD.t1551 557.608
R5898 VDD.t1221 VDD.t871 556.306
R5899 VDD.t1763 VDD.t1203 556.306
R5900 VDD.t919 VDD.t1207 556.306
R5901 VDD.t1353 VDD.t1195 556.306
R5902 VDD.t845 VDD.t1223 556.306
R5903 VDD.t1005 VDD.t1209 556.306
R5904 VDD.t1433 VDD.t1213 556.306
R5905 VDD.t635 VDD.t1199 556.306
R5906 VDD.t2278 VDD.t1215 544.894
R5907 VDD.t1531 VDD.t1217 544.894
R5908 VDD.t2270 VDD.t1201 544.894
R5909 VDD.t1288 VDD.t1205 544.894
R5910 VDD.t1504 VDD.t1193 544.894
R5911 VDD.t1814 VDD.t1197 544.894
R5912 VDD.t334 VDD.t1219 544.894
R5913 VDD.t2165 VDD.t1211 518.181
R5914 VDD.t1832 VDD.t1154 509.926
R5915 VDD.t431 VDD.t1124 509.926
R5916 VDD.t1787 VDD.t1130 509.926
R5917 VDD.t1981 VDD.t1104 509.926
R5918 VDD.t1580 VDD.t1134 509.926
R5919 VDD.t30 VDD.t1106 509.926
R5920 VDD.t1072 VDD.t1110 509.926
R5921 VDD.t1399 VDD.t1132 509.926
R5922 VDD.t4 VDD.t1116 509.926
R5923 VDD.t1060 VDD.t1136 509.926
R5924 VDD.t336 VDD.t1158 509.926
R5925 VDD.t1456 VDD.t1112 509.926
R5926 VDD.t752 VDD.t1164 509.926
R5927 VDD.t2109 VDD.t1120 509.926
R5928 VDD.t1710 VDD.t1128 509.926
R5929 VDD.t1675 VDD.t1152 509.926
R5930 VDD.t619 VDD.t1146 499.448
R5931 VDD.t1235 VDD.t1114 499.448
R5932 VDD.t1789 VDD.t1148 499.448
R5933 VDD.t1797 VDD.t1156 499.448
R5934 VDD.t571 VDD.t1126 499.448
R5935 VDD.t512 VDD.t1162 499.448
R5936 VDD.t427 VDD.t1118 499.448
R5937 VDD.t1172 VDD.t1138 499.448
R5938 VDD.t1176 VDD.t1160 499.448
R5939 VDD.t1319 VDD.t1142 499.448
R5940 VDD.t2194 VDD.t1166 499.448
R5941 VDD.t741 VDD.t1122 499.448
R5942 VDD.t326 VDD.t1140 499.448
R5943 VDD.t2258 VDD.t1108 499.448
R5944 VDD.t1698 VDD.t1144 499.448
R5945 VDD.t1182 VDD.t1150 499.448
R5946 VDD.t2056 VDD.t2063 475
R5947 VDD.t2022 VDD.t2028 475
R5948 VDD.t2043 VDD.t2026 475
R5949 VDD.t2083 VDD.t2089 475
R5950 VDD.t2025 VDD.t2034 475
R5951 VDD.t2088 VDD.t2020 475
R5952 VDD.t2087 VDD.t2018 475
R5953 VDD.t2075 VDD.t2081 475
R5954 VDD.t2017 VDD.t2023 475
R5955 VDD.t2055 VDD.t2061 475
R5956 VDD.t2080 VDD.t2085 475
R5957 VDD.t2042 VDD.t2049 475
R5958 VDD.t2084 VDD.t2015 475
R5959 VDD.t2048 VDD.t2053 475
R5960 VDD.t2074 VDD.t2078 475
R5961 VDD.t2065 VDD.t2068 475
R5962 VDD.n588 VDD.t2032 465.104
R5963 VDD.n660 VDD.t2046 465.104
R5964 VDD.n732 VDD.t2011 465.104
R5965 VDD.n804 VDD.t2038 465.104
R5966 VDD.n876 VDD.t2072 465.104
R5967 VDD.n948 VDD.t2040 465.104
R5968 VDD.n1020 VDD.t2059 465.104
R5969 VDD.n1092 VDD.t2030 465.104
R5970 VDD.n1164 VDD.t2066 465.104
R5971 VDD.n1236 VDD.t2036 465.104
R5972 VDD.n1308 VDD.t2051 465.104
R5973 VDD.n1380 VDD.t2070 465.104
R5974 VDD.n1452 VDD.t2057 465.104
R5975 VDD.n1524 VDD.t2076 465.104
R5976 VDD.n1596 VDD.t2044 465.104
R5977 VDD.n1607 VDD.t2013 465.104
R5978 VDD.n595 VDD.t2033 416.315
R5979 VDD.n739 VDD.t2012 416.315
R5980 VDD.n811 VDD.t2039 416.315
R5981 VDD.n883 VDD.t2073 416.315
R5982 VDD.n955 VDD.t2041 416.315
R5983 VDD.n1027 VDD.t2060 416.315
R5984 VDD.n1099 VDD.t2031 416.315
R5985 VDD.n1171 VDD.t2067 416.315
R5986 VDD.n1243 VDD.t2037 416.315
R5987 VDD.n1315 VDD.t2052 416.315
R5988 VDD.n1387 VDD.t2071 416.315
R5989 VDD.n1459 VDD.t2058 416.315
R5990 VDD.n1531 VDD.t2077 416.315
R5991 VDD.n1603 VDD.t2045 416.315
R5992 VDD.n1606 VDD.t2014 416.315
R5993 VDD.n667 VDD.t2047 416.315
R5994 VDD.n595 VDD.t2064 416.142
R5995 VDD.n739 VDD.t2027 416.142
R5996 VDD.n811 VDD.t2090 416.142
R5997 VDD.n883 VDD.t2035 416.142
R5998 VDD.n955 VDD.t2021 416.142
R5999 VDD.n1027 VDD.t2019 416.142
R6000 VDD.n1099 VDD.t2082 416.142
R6001 VDD.n1171 VDD.t2024 416.142
R6002 VDD.n1243 VDD.t2062 416.142
R6003 VDD.n1315 VDD.t2086 416.142
R6004 VDD.n1387 VDD.t2050 416.142
R6005 VDD.n1459 VDD.t2016 416.142
R6006 VDD.n1531 VDD.t2054 416.142
R6007 VDD.n1603 VDD.t2079 416.142
R6008 VDD.n1606 VDD.t2069 416.142
R6009 VDD.n667 VDD.t2029 416.142
R6010 VDD.t1307 VDD.t184 298.189
R6011 VDD.t1553 VDD.t236 298.189
R6012 VDD.t1596 VDD.t182 298.189
R6013 VDD.t1447 VDD.t232 298.189
R6014 VDD.t2095 VDD.t294 298.189
R6015 VDD.t419 VDD.t126 298.189
R6016 VDD.t1535 VDD.t142 298.189
R6017 VDD.t76 VDD.t190 298.189
R6018 VDD.t1653 VDD.t112 298.189
R6019 VDD.t663 VDD.t156 298.189
R6020 VDD.t397 VDD.t238 298.189
R6021 VDD.t723 VDD.t265 298.189
R6022 VDD.t1444 VDD.t154 298.189
R6023 VDD.t1997 VDD.t200 298.189
R6024 VDD.t849 VDD.t292 298.189
R6025 VDD.t1096 VDD.t122 298.189
R6026 VDD.t1749 VDD.t180 298.189
R6027 VDD.t997 VDD.t230 298.189
R6028 VDD.t366 VDD.t259 298.189
R6029 VDD.t1977 VDD.t286 298.189
R6030 VDD.t1727 VDD.t162 298.189
R6031 VDD.t699 VDD.t206 298.189
R6032 VDD.t1018 VDD.t178 298.189
R6033 VDD.t1082 VDD.t228 298.189
R6034 VDD.t1567 VDD.t192 298.189
R6035 VDD.t1315 VDD.t240 298.189
R6036 VDD.t2260 VDD.t170 298.189
R6037 VDD.t1834 VDD.t216 298.189
R6038 VDD.t1371 VDD.t221 298.189
R6039 VDD.t1290 VDD.t254 298.189
R6040 VDD.t861 VDD.t164 298.189
R6041 VDD.t1335 VDD.t209 298.189
R6042 VDD.t274 VDD.t1419 292.454
R6043 VDD.t304 VDD.t915 292.454
R6044 VDD.t270 VDD.t1070 292.454
R6045 VDD.t302 VDD.t1449 292.454
R6046 VDD.t124 VDD.t543 292.454
R6047 VDD.t166 VDD.t1639 292.454
R6048 VDD.t277 VDD.t1537 292.454
R6049 VDD.t86 VDD.t1068 292.454
R6050 VDD.t261 VDD.t1381 292.454
R6051 VDD.t288 VDD.t665 292.454
R6052 VDD.t132 VDD.t1466 292.454
R6053 VDD.t174 VDD.t719 292.454
R6054 VDD.t281 VDD.t811 292.454
R6055 VDD.t90 VDD.t1180 292.454
R6056 VDD.t223 VDD.t893 292.454
R6057 VDD.t257 VDD.t1619 292.454
R6058 VDD.t116 VDD.t1549 292.454
R6059 VDD.t160 VDD.t789 292.454
R6060 VDD.t202 VDD.t1253 292.454
R6061 VDD.t245 VDD.t1979 292.454
R6062 VDD.t283 VDD.t1510 292.454
R6063 VDD.t102 VDD.t348 292.454
R6064 VDD.t298 VDD.t551 292.454
R6065 VDD.t130 VDD.t1850 292.454
R6066 VDD.t148 VDD.t1451 292.454
R6067 VDD.t196 VDD.t1317 292.454
R6068 VDD.t108 VDD.t2105 292.454
R6069 VDD.t152 VDD.t847 292.454
R6070 VDD.t308 VDD.t1441 292.454
R6071 VDD.t134 VDD.t1294 292.454
R6072 VDD.t267 VDD.t1030 292.454
R6073 VDD.t296 VDD.t1337 292.454
R6074 VDD.n1541 VDD.t1763 282.432
R6075 VDD.n1397 VDD.t919 282.432
R6076 VDD.n1253 VDD.t1353 282.432
R6077 VDD.n1109 VDD.t845 282.432
R6078 VDD.n965 VDD.t1005 282.432
R6079 VDD.n821 VDD.t1433 282.432
R6080 VDD.n677 VDD.t635 282.432
R6081 VDD.n1541 VDD.t2278 256.756
R6082 VDD.n1397 VDD.t1531 256.756
R6083 VDD.n1253 VDD.t2270 256.756
R6084 VDD.n1109 VDD.t1288 256.756
R6085 VDD.n965 VDD.t1504 256.756
R6086 VDD.n821 VDD.t1814 256.756
R6087 VDD.n677 VDD.t334 256.756
R6088 VDD.n539 VDD.t2166 250.672
R6089 VDD.n604 VDD.t636 250.092
R6090 VDD.n679 VDD.t1242 250.092
R6091 VDD.n751 VDD.t1434 250.092
R6092 VDD.n823 VDD.t626 250.092
R6093 VDD.n895 VDD.t1006 250.092
R6094 VDD.n967 VDD.t1857 250.092
R6095 VDD.n1039 VDD.t846 250.092
R6096 VDD.n1111 VDD.t1766 250.092
R6097 VDD.n1183 VDD.t1354 250.092
R6098 VDD.n1255 VDD.t860 250.092
R6099 VDD.n1327 VDD.t920 250.092
R6100 VDD.n1399 VDD.t1053 250.092
R6101 VDD.n1471 VDD.t1764 250.092
R6102 VDD.n1543 VDD.t2287 250.092
R6103 VDD.n1623 VDD.t872 250.092
R6104 VDD.n678 VDD.t335 244.267
R6105 VDD.n750 VDD.t1252 244.267
R6106 VDD.n822 VDD.t1815 244.267
R6107 VDD.n894 VDD.t511 244.267
R6108 VDD.n966 VDD.t1505 244.267
R6109 VDD.n1038 VDD.t874 244.267
R6110 VDD.n1110 VDD.t1289 244.267
R6111 VDD.n1182 VDD.t498 244.267
R6112 VDD.n1254 VDD.t2271 244.267
R6113 VDD.n1326 VDD.t804 244.267
R6114 VDD.n1398 VDD.t1532 244.267
R6115 VDD.n1470 VDD.t2092 244.267
R6116 VDD.n1542 VDD.t2279 244.267
R6117 VDD.n603 VDD.t638 244.267
R6118 VDD.n1622 VDD.t556 243.928
R6119 VDD.n538 VDD.t1004 241.449
R6120 VDD.n1622 VDD.n1621 229.589
R6121 VDD.n734 VDD.n733 229.55
R6122 VDD.n806 VDD.n805 229.55
R6123 VDD.n878 VDD.n877 229.55
R6124 VDD.n950 VDD.n949 229.55
R6125 VDD.n1022 VDD.n1021 229.55
R6126 VDD.n1094 VDD.n1093 229.55
R6127 VDD.n1166 VDD.n1165 229.55
R6128 VDD.n1238 VDD.n1237 229.55
R6129 VDD.n1310 VDD.n1309 229.55
R6130 VDD.n1382 VDD.n1381 229.55
R6131 VDD.n1454 VDD.n1453 229.55
R6132 VDD.n1526 VDD.n1525 229.55
R6133 VDD.n1598 VDD.n1597 229.55
R6134 VDD.n662 VDD.n661 229.55
R6135 VDD.n701 VDD.n700 229.55
R6136 VDD.n719 VDD.n718 229.55
R6137 VDD.n672 VDD.n671 229.55
R6138 VDD.n773 VDD.n772 229.55
R6139 VDD.n791 VDD.n790 229.55
R6140 VDD.n744 VDD.n743 229.55
R6141 VDD.n845 VDD.n844 229.55
R6142 VDD.n863 VDD.n862 229.55
R6143 VDD.n816 VDD.n815 229.55
R6144 VDD.n917 VDD.n916 229.55
R6145 VDD.n935 VDD.n934 229.55
R6146 VDD.n888 VDD.n887 229.55
R6147 VDD.n989 VDD.n988 229.55
R6148 VDD.n1007 VDD.n1006 229.55
R6149 VDD.n960 VDD.n959 229.55
R6150 VDD.n1061 VDD.n1060 229.55
R6151 VDD.n1079 VDD.n1078 229.55
R6152 VDD.n1032 VDD.n1031 229.55
R6153 VDD.n1133 VDD.n1132 229.55
R6154 VDD.n1151 VDD.n1150 229.55
R6155 VDD.n1104 VDD.n1103 229.55
R6156 VDD.n1205 VDD.n1204 229.55
R6157 VDD.n1223 VDD.n1222 229.55
R6158 VDD.n1176 VDD.n1175 229.55
R6159 VDD.n1277 VDD.n1276 229.55
R6160 VDD.n1295 VDD.n1294 229.55
R6161 VDD.n1248 VDD.n1247 229.55
R6162 VDD.n1349 VDD.n1348 229.55
R6163 VDD.n1367 VDD.n1366 229.55
R6164 VDD.n1320 VDD.n1319 229.55
R6165 VDD.n1421 VDD.n1420 229.55
R6166 VDD.n1439 VDD.n1438 229.55
R6167 VDD.n1392 VDD.n1391 229.55
R6168 VDD.n1493 VDD.n1492 229.55
R6169 VDD.n1511 VDD.n1510 229.55
R6170 VDD.n1464 VDD.n1463 229.55
R6171 VDD.n1565 VDD.n1564 229.55
R6172 VDD.n1583 VDD.n1582 229.55
R6173 VDD.n1536 VDD.n1535 229.55
R6174 VDD.n1609 VDD.n1608 229.55
R6175 VDD.n1611 VDD.n1610 229.55
R6176 VDD.n1613 VDD.n1612 229.55
R6177 VDD.n1616 VDD.n1615 229.55
R6178 VDD.n528 VDD.n527 229.55
R6179 VDD.n530 VDD.n529 229.55
R6180 VDD.n533 VDD.n532 229.55
R6181 VDD.n615 VDD.n614 229.55
R6182 VDD.n629 VDD.n628 229.55
R6183 VDD.n647 VDD.n646 229.55
R6184 VDD.n590 VDD.n589 229.55
R6185 VDD.n678 VDD.n677 229.423
R6186 VDD.n750 VDD.n749 229.423
R6187 VDD.n822 VDD.n821 229.423
R6188 VDD.n894 VDD.n893 229.423
R6189 VDD.n966 VDD.n965 229.423
R6190 VDD.n1038 VDD.n1037 229.423
R6191 VDD.n1110 VDD.n1109 229.423
R6192 VDD.n1182 VDD.n1181 229.423
R6193 VDD.n1254 VDD.n1253 229.423
R6194 VDD.n1326 VDD.n1325 229.423
R6195 VDD.n1398 VDD.n1397 229.423
R6196 VDD.n1470 VDD.n1469 229.423
R6197 VDD.n1542 VDD.n1541 229.423
R6198 VDD.n99 VDD.t277 189.546
R6199 VDD.n131 VDD.t261 189.546
R6200 VDD.n163 VDD.t132 189.546
R6201 VDD.n195 VDD.t281 189.546
R6202 VDD.n227 VDD.t223 189.546
R6203 VDD.n259 VDD.t116 189.546
R6204 VDD.n291 VDD.t202 189.546
R6205 VDD.n323 VDD.t283 189.546
R6206 VDD.n355 VDD.t298 189.546
R6207 VDD.n387 VDD.t148 189.546
R6208 VDD.n419 VDD.t108 189.546
R6209 VDD.n451 VDD.t308 189.546
R6210 VDD.n483 VDD.t267 189.546
R6211 VDD.n3 VDD.t274 187.635
R6212 VDD.n35 VDD.t270 187.635
R6213 VDD.n67 VDD.t124 187.635
R6214 VDD.t1419 VDD.t1307 185.412
R6215 VDD.t915 VDD.t1553 185.412
R6216 VDD.t1070 VDD.t1596 185.412
R6217 VDD.t1449 VDD.t1447 185.412
R6218 VDD.t543 VDD.t2095 185.412
R6219 VDD.t1639 VDD.t419 185.412
R6220 VDD.t1381 VDD.t1653 185.412
R6221 VDD.t665 VDD.t663 185.412
R6222 VDD.t1466 VDD.t397 185.412
R6223 VDD.t719 VDD.t723 185.412
R6224 VDD.t811 VDD.t1444 185.412
R6225 VDD.t1180 VDD.t1997 185.412
R6226 VDD.t893 VDD.t849 185.412
R6227 VDD.t1619 VDD.t1096 185.412
R6228 VDD.t1549 VDD.t1749 185.412
R6229 VDD.t789 VDD.t997 185.412
R6230 VDD.t1253 VDD.t366 185.412
R6231 VDD.t1979 VDD.t1977 185.412
R6232 VDD.t1510 VDD.t1727 185.412
R6233 VDD.t348 VDD.t699 185.412
R6234 VDD.t551 VDD.t1018 185.412
R6235 VDD.t1850 VDD.t1082 185.412
R6236 VDD.t1451 VDD.t1567 185.412
R6237 VDD.t1317 VDD.t1315 185.412
R6238 VDD.t2105 VDD.t2260 185.412
R6239 VDD.t847 VDD.t1834 185.412
R6240 VDD.t1441 VDD.t1371 185.412
R6241 VDD.t1294 VDD.t1290 185.412
R6242 VDD.t1030 VDD.t861 185.412
R6243 VDD.t1337 VDD.t1335 185.412
R6244 VDD.n602 VDD.n601 185
R6245 VDD.t1537 VDD.t1535 183.501
R6246 VDD.t1068 VDD.t76 183.501
R6247 VDD.n109 VDD.t86 179.945
R6248 VDD.n141 VDD.t288 179.945
R6249 VDD.n173 VDD.t174 179.945
R6250 VDD.n205 VDD.t90 179.945
R6251 VDD.n237 VDD.t257 179.945
R6252 VDD.n269 VDD.t160 179.945
R6253 VDD.n301 VDD.t245 179.945
R6254 VDD.n333 VDD.t102 179.945
R6255 VDD.n365 VDD.t130 179.945
R6256 VDD.n397 VDD.t196 179.945
R6257 VDD.n429 VDD.t152 179.945
R6258 VDD.n461 VDD.t134 179.945
R6259 VDD.n493 VDD.t296 179.945
R6260 VDD.n13 VDD.t304 178.033
R6261 VDD.n45 VDD.t302 178.033
R6262 VDD.n77 VDD.t166 178.033
R6263 VDD.n531 VDD.t1832 171.139
R6264 VDD.n613 VDD.t431 171.139
R6265 VDD.n670 VDD.t1787 171.139
R6266 VDD.n742 VDD.t1981 171.139
R6267 VDD.n814 VDD.t1580 171.139
R6268 VDD.n886 VDD.t30 171.139
R6269 VDD.n958 VDD.t1072 171.139
R6270 VDD.n1030 VDD.t1399 171.139
R6271 VDD.n1102 VDD.t4 171.139
R6272 VDD.n1174 VDD.t1060 171.139
R6273 VDD.n1246 VDD.t336 171.139
R6274 VDD.n1318 VDD.t1456 171.139
R6275 VDD.n1390 VDD.t752 171.139
R6276 VDD.n1462 VDD.t2109 171.139
R6277 VDD.n1534 VDD.t1710 171.139
R6278 VDD.n1614 VDD.t1675 171.139
R6279 VDD.n531 VDD.t619 167.647
R6280 VDD.n613 VDD.t1235 167.647
R6281 VDD.n670 VDD.t1789 167.647
R6282 VDD.n742 VDD.t1797 167.647
R6283 VDD.n814 VDD.t571 167.647
R6284 VDD.n886 VDD.t512 167.647
R6285 VDD.n958 VDD.t427 167.647
R6286 VDD.n1030 VDD.t1172 167.647
R6287 VDD.n1102 VDD.t1176 167.647
R6288 VDD.n1174 VDD.t1319 167.647
R6289 VDD.n1246 VDD.t2194 167.647
R6290 VDD.n1318 VDD.t741 167.647
R6291 VDD.n1390 VDD.t326 167.647
R6292 VDD.n1462 VDD.t2258 167.647
R6293 VDD.n1534 VDD.t1698 167.647
R6294 VDD.n1614 VDD.t1182 167.647
R6295 VDD.n1 VDD.t1308 156.041
R6296 VDD.n5 VDD.t394 156.041
R6297 VDD.n32 VDD.t1597 156.041
R6298 VDD.n38 VDD.t1045 156.041
R6299 VDD.n65 VDD.t2096 156.041
R6300 VDD.n69 VDD.t2276 156.041
R6301 VDD.n96 VDD.t1536 156.041
R6302 VDD.n101 VDD.t1530 156.041
R6303 VDD.n128 VDD.t1654 156.041
R6304 VDD.n133 VDD.t1446 156.041
R6305 VDD.n161 VDD.t398 156.041
R6306 VDD.n166 VDD.t1646 156.041
R6307 VDD.n192 VDD.t1445 156.041
R6308 VDD.n197 VDD.t1009 156.041
R6309 VDD.n224 VDD.t850 156.041
R6310 VDD.n229 VDD.t1263 156.041
R6311 VDD.n256 VDD.t1750 156.041
R6312 VDD.n262 VDD.t1455 156.041
R6313 VDD.n288 VDD.t367 156.041
R6314 VDD.n293 VDD.t624 156.041
R6315 VDD.n320 VDD.t1728 156.041
R6316 VDD.n326 VDD.t73 156.041
R6317 VDD.n353 VDD.t1019 156.041
R6318 VDD.n357 VDD.t2245 156.041
R6319 VDD.n385 VDD.t1568 156.041
R6320 VDD.n390 VDD.t1509 156.041
R6321 VDD.n417 VDD.t2261 156.041
R6322 VDD.n421 VDD.t61 156.041
R6323 VDD.n448 VDD.t1372 156.041
R6324 VDD.n454 VDD.t1807 156.041
R6325 VDD.n481 VDD.t862 156.041
R6326 VDD.n485 VDD.t1037 156.041
R6327 VDD.n26 VDD.t363 155.985
R6328 VDD.n11 VDD.t1554 155.985
R6329 VDD.n58 VDD.t1416 155.985
R6330 VDD.n43 VDD.t1448 155.985
R6331 VDD.n90 VDD.t1591 155.985
R6332 VDD.n75 VDD.t420 155.985
R6333 VDD.n122 VDD.t878 155.985
R6334 VDD.n107 VDD.t77 155.985
R6335 VDD.n154 VDD.t1271 155.985
R6336 VDD.n139 VDD.t664 155.985
R6337 VDD.n186 VDD.t798 155.985
R6338 VDD.n171 VDD.t724 155.985
R6339 VDD.n218 VDD.t402 155.985
R6340 VDD.n203 VDD.t1998 155.985
R6341 VDD.n250 VDD.t1085 155.985
R6342 VDD.n235 VDD.t1097 155.985
R6343 VDD.n282 VDD.t980 155.985
R6344 VDD.n267 VDD.t998 155.985
R6345 VDD.n314 VDD.t1677 155.985
R6346 VDD.n299 VDD.t1978 155.985
R6347 VDD.n346 VDD.t518 155.985
R6348 VDD.n331 VDD.t700 155.985
R6349 VDD.n378 VDD.t1656 155.985
R6350 VDD.n363 VDD.t1083 155.985
R6351 VDD.n410 VDD.t1868 155.985
R6352 VDD.n395 VDD.t1316 155.985
R6353 VDD.n442 VDD.t1610 155.985
R6354 VDD.n427 VDD.t1835 155.985
R6355 VDD.n474 VDD.t566 155.985
R6356 VDD.n459 VDD.t1291 155.985
R6357 VDD.n506 VDD.t2183 155.985
R6358 VDD.n491 VDD.t1336 155.985
R6359 VDD.t362 VDD.t104 155.508
R6360 VDD.t1044 VDD.t98 155.508
R6361 VDD.t1590 VDD.t144 155.508
R6362 VDD.t877 VDD.t211 155.508
R6363 VDD.t1270 VDD.t172 155.508
R6364 VDD.t797 VDD.t150 155.508
R6365 VDD.t401 VDD.t219 155.508
R6366 VDD.t1084 VDD.t140 155.508
R6367 VDD.t979 VDD.t96 155.508
R6368 VDD.t623 VDD.t186 155.508
R6369 VDD.t72 VDD.t226 155.508
R6370 VDD.t1655 VDD.t94 155.508
R6371 VDD.t1508 VDD.t110 155.508
R6372 VDD.t60 VDD.t88 155.508
R6373 VDD.t565 VDD.t136 155.508
R6374 VDD.t1036 VDD.t234 155.508
R6375 VDD.n1 VDD.t1420 155.288
R6376 VDD.n5 VDD.t365 155.288
R6377 VDD.n32 VDD.t1071 155.288
R6378 VDD.n38 VDD.t1403 155.288
R6379 VDD.n65 VDD.t544 155.288
R6380 VDD.n69 VDD.t2277 155.288
R6381 VDD.n96 VDD.t1538 155.288
R6382 VDD.n101 VDD.t682 155.288
R6383 VDD.n128 VDD.t1382 155.288
R6384 VDD.n133 VDD.t828 155.288
R6385 VDD.n161 VDD.t1467 155.288
R6386 VDD.n166 VDD.t1645 155.288
R6387 VDD.n192 VDD.t812 155.288
R6388 VDD.n197 VDD.t1055 155.288
R6389 VDD.n224 VDD.t894 155.288
R6390 VDD.n229 VDD.t1228 155.288
R6391 VDD.n256 VDD.t1550 155.288
R6392 VDD.n262 VDD.t472 155.288
R6393 VDD.n288 VDD.t1254 155.288
R6394 VDD.n293 VDD.t1712 155.288
R6395 VDD.n320 VDD.t1511 155.288
R6396 VDD.n326 VDD.t23 155.288
R6397 VDD.n353 VDD.t552 155.288
R6398 VDD.n357 VDD.t2230 155.288
R6399 VDD.n385 VDD.t1452 155.288
R6400 VDD.n390 VDD.t1277 155.288
R6401 VDD.n417 VDD.t2106 155.288
R6402 VDD.n421 VDD.t33 155.288
R6403 VDD.n448 VDD.t1442 155.288
R6404 VDD.n454 VDD.t1601 155.288
R6405 VDD.n481 VDD.t1031 155.288
R6406 VDD.n485 VDD.t1088 155.288
R6407 VDD.n26 VDD.t788 155.232
R6408 VDD.n11 VDD.t916 155.232
R6409 VDD.n58 VDD.t426 155.232
R6410 VDD.n43 VDD.t1450 155.232
R6411 VDD.n90 VDD.t1776 155.232
R6412 VDD.n75 VDD.t1640 155.232
R6413 VDD.n122 VDD.t743 155.232
R6414 VDD.n107 VDD.t1069 155.232
R6415 VDD.n154 VDD.t1600 155.232
R6416 VDD.n139 VDD.t666 155.232
R6417 VDD.n186 VDD.t747 155.232
R6418 VDD.n171 VDD.t720 155.232
R6419 VDD.n218 VDD.t1192 155.232
R6420 VDD.n203 VDD.t1181 155.232
R6421 VDD.n250 VDD.t1571 155.232
R6422 VDD.n235 VDD.t1620 155.232
R6423 VDD.n282 VDD.t1089 155.232
R6424 VDD.n267 VDD.t790 155.232
R6425 VDD.n314 VDD.t1674 155.232
R6426 VDD.n299 VDD.t1980 155.232
R6427 VDD.n346 VDD.t1443 155.232
R6428 VDD.n331 VDD.t349 155.232
R6429 VDD.n378 VDD.t1430 155.232
R6430 VDD.n363 VDD.t1851 155.232
R6431 VDD.n410 VDD.t1296 155.232
R6432 VDD.n395 VDD.t1318 155.232
R6433 VDD.n442 VDD.t509 155.232
R6434 VDD.n427 VDD.t848 155.232
R6435 VDD.n474 VDD.t1238 155.232
R6436 VDD.n459 VDD.t1295 155.232
R6437 VDD.n506 VDD.t19 155.232
R6438 VDD.n491 VDD.t1338 155.232
R6439 VDD.t106 VDD.t364 152.518
R6440 VDD.t100 VDD.t425 152.518
R6441 VDD.t188 VDD.t1775 152.518
R6442 VDD.t114 VDD.t681 152.518
R6443 VDD.t194 VDD.t827 152.518
R6444 VDD.t198 VDD.t746 152.518
R6445 VDD.t118 VDD.t1054 152.518
R6446 VDD.t138 VDD.t1227 152.518
R6447 VDD.t176 VDD.t471 152.518
R6448 VDD.t120 VDD.t1673 152.518
R6449 VDD.t128 VDD.t22 152.518
R6450 VDD.t146 VDD.t1429 152.518
R6451 VDD.t214 VDD.t1276 152.518
R6452 VDD.t168 VDD.t32 152.518
R6453 VDD.t158 VDD.t1237 152.518
R6454 VDD.t92 VDD.t18 152.518
R6455 VDD.n0 VDD.t185 144.383
R6456 VDD.n7 VDD.t105 144.383
R6457 VDD.n34 VDD.t183 144.383
R6458 VDD.n37 VDD.t99 144.383
R6459 VDD.n64 VDD.t295 144.383
R6460 VDD.n71 VDD.t244 144.383
R6461 VDD.n98 VDD.t143 144.383
R6462 VDD.n103 VDD.t285 144.383
R6463 VDD.n130 VDD.t113 144.383
R6464 VDD.n135 VDD.t264 144.383
R6465 VDD.n160 VDD.t239 144.383
R6466 VDD.n165 VDD.t151 144.383
R6467 VDD.n194 VDD.t155 144.383
R6468 VDD.n199 VDD.t291 144.383
R6469 VDD.n226 VDD.t293 144.383
R6470 VDD.n231 VDD.t243 144.383
R6471 VDD.n258 VDD.t181 144.383
R6472 VDD.n261 VDD.t97 144.383
R6473 VDD.n290 VDD.t260 144.383
R6474 VDD.n295 VDD.t187 144.383
R6475 VDD.n322 VDD.t163 144.383
R6476 VDD.n325 VDD.t300 144.383
R6477 VDD.n352 VDD.t179 144.383
R6478 VDD.n359 VDD.t95 144.383
R6479 VDD.n384 VDD.t193 144.383
R6480 VDD.n389 VDD.t111 144.383
R6481 VDD.n416 VDD.t171 144.383
R6482 VDD.n423 VDD.t89 144.383
R6483 VDD.n450 VDD.t222 144.383
R6484 VDD.n453 VDD.t137 144.383
R6485 VDD.n480 VDD.t165 144.383
R6486 VDD.n487 VDD.t301 144.383
R6487 VDD.n25 VDD.t251 144.291
R6488 VDD.n10 VDD.t237 144.291
R6489 VDD.n57 VDD.t250 144.291
R6490 VDD.n42 VDD.t233 144.291
R6491 VDD.n89 VDD.t145 144.291
R6492 VDD.n74 VDD.t127 144.291
R6493 VDD.n121 VDD.t212 144.291
R6494 VDD.n106 VDD.t191 144.291
R6495 VDD.n153 VDD.t173 144.291
R6496 VDD.n138 VDD.t157 144.291
R6497 VDD.n185 VDD.t280 144.291
R6498 VDD.n170 VDD.t266 144.291
R6499 VDD.n217 VDD.t220 144.291
R6500 VDD.n202 VDD.t201 144.291
R6501 VDD.n249 VDD.t141 144.291
R6502 VDD.n234 VDD.t123 144.291
R6503 VDD.n281 VDD.t249 144.291
R6504 VDD.n266 VDD.t231 144.291
R6505 VDD.n313 VDD.t306 144.291
R6506 VDD.n298 VDD.t287 144.291
R6507 VDD.n345 VDD.t227 144.291
R6508 VDD.n330 VDD.t207 144.291
R6509 VDD.n377 VDD.t248 144.291
R6510 VDD.n362 VDD.t229 144.291
R6511 VDD.n409 VDD.t252 144.291
R6512 VDD.n394 VDD.t241 144.291
R6513 VDD.n441 VDD.t242 144.291
R6514 VDD.n426 VDD.t217 144.291
R6515 VDD.n473 VDD.t272 144.291
R6516 VDD.n458 VDD.t255 144.291
R6517 VDD.n505 VDD.t235 144.291
R6518 VDD.n490 VDD.t210 144.291
R6519 VDD.n3 VDD.t275 142.941
R6520 VDD.n8 VDD.t208 142.941
R6521 VDD.n35 VDD.t271 142.941
R6522 VDD.n40 VDD.t205 142.941
R6523 VDD.n67 VDD.t125 142.941
R6524 VDD.n72 VDD.t276 142.941
R6525 VDD.n99 VDD.t278 142.941
R6526 VDD.n104 VDD.t213 142.941
R6527 VDD.n131 VDD.t262 142.941
R6528 VDD.n136 VDD.t195 142.941
R6529 VDD.n163 VDD.t133 142.941
R6530 VDD.n168 VDD.t279 142.941
R6531 VDD.n195 VDD.t282 142.941
R6532 VDD.n200 VDD.t218 142.941
R6533 VDD.n227 VDD.t224 142.941
R6534 VDD.n232 VDD.t139 142.941
R6535 VDD.n259 VDD.t117 142.941
R6536 VDD.n264 VDD.t269 142.941
R6537 VDD.n291 VDD.t203 142.941
R6538 VDD.n296 VDD.t121 142.941
R6539 VDD.n323 VDD.t284 142.941
R6540 VDD.n328 VDD.t225 142.941
R6541 VDD.n355 VDD.t299 142.941
R6542 VDD.n360 VDD.t247 142.941
R6543 VDD.n387 VDD.t149 142.941
R6544 VDD.n392 VDD.t290 142.941
R6545 VDD.n419 VDD.t109 142.941
R6546 VDD.n424 VDD.t263 142.941
R6547 VDD.n451 VDD.t309 142.941
R6548 VDD.n456 VDD.t253 142.941
R6549 VDD.n483 VDD.t268 142.941
R6550 VDD.n488 VDD.t204 142.941
R6551 VDD.n23 VDD.t107 142.93
R6552 VDD.n13 VDD.t305 142.93
R6553 VDD.n55 VDD.t101 142.93
R6554 VDD.n45 VDD.t303 142.93
R6555 VDD.n87 VDD.t189 142.93
R6556 VDD.n77 VDD.t167 142.93
R6557 VDD.n119 VDD.t115 142.93
R6558 VDD.n109 VDD.t87 142.93
R6559 VDD.n151 VDD.t307 142.93
R6560 VDD.n141 VDD.t289 142.93
R6561 VDD.n183 VDD.t199 142.93
R6562 VDD.n173 VDD.t175 142.93
R6563 VDD.n215 VDD.t119 142.93
R6564 VDD.n205 VDD.t91 142.93
R6565 VDD.n247 VDD.t273 142.93
R6566 VDD.n237 VDD.t258 142.93
R6567 VDD.n279 VDD.t177 142.93
R6568 VDD.n269 VDD.t161 142.93
R6569 VDD.n311 VDD.t256 142.93
R6570 VDD.n301 VDD.t246 142.93
R6571 VDD.n343 VDD.t129 142.93
R6572 VDD.n333 VDD.t103 142.93
R6573 VDD.n375 VDD.t147 142.93
R6574 VDD.n365 VDD.t131 142.93
R6575 VDD.n407 VDD.t215 142.93
R6576 VDD.n397 VDD.t197 142.93
R6577 VDD.n439 VDD.t169 142.93
R6578 VDD.n429 VDD.t153 142.93
R6579 VDD.n471 VDD.t159 142.93
R6580 VDD.n461 VDD.t135 142.93
R6581 VDD.n503 VDD.t93 142.93
R6582 VDD.n493 VDD.t297 142.93
R6583 VDD.n690 VDD.t2263 102.87
R6584 VDD.n692 VDD.t794 102.87
R6585 VDD.n694 VDD.t974 102.87
R6586 VDD.n696 VDD.t2205 102.87
R6587 VDD.n698 VDD.t968 102.87
R6588 VDD.n704 VDD.t454 102.87
R6589 VDD.n706 VDD.t938 102.87
R6590 VDD.n708 VDD.t1853 102.87
R6591 VDD.n710 VDD.t1644 102.87
R6592 VDD.n712 VDD.t1023 102.87
R6593 VDD.n714 VDD.t1884 102.87
R6594 VDD.n716 VDD.t1507 102.87
R6595 VDD.n722 VDD.t474 102.87
R6596 VDD.n724 VDD.t1966 102.87
R6597 VDD.n726 VDD.t1593 102.87
R6598 VDD.n728 VDD.t29 102.87
R6599 VDD.n730 VDD.t978 102.87
R6600 VDD.n737 VDD.t492 102.87
R6601 VDD.n686 VDD.t767 102.87
R6602 VDD.n684 VDD.t785 102.87
R6603 VDD.n762 VDD.t2160 102.87
R6604 VDD.n764 VDD.t775 102.87
R6605 VDD.n766 VDD.t63 102.87
R6606 VDD.n768 VDD.t728 102.87
R6607 VDD.n770 VDD.t2142 102.87
R6608 VDD.n776 VDD.t554 102.87
R6609 VDD.n778 VDD.t438 102.87
R6610 VDD.n780 VDD.t781 102.87
R6611 VDD.n782 VDD.t1169 102.87
R6612 VDD.n784 VDD.t2225 102.87
R6613 VDD.n786 VDD.t2176 102.87
R6614 VDD.n788 VDD.t884 102.87
R6615 VDD.n794 VDD.t1185 102.87
R6616 VDD.n796 VDD.t1388 102.87
R6617 VDD.n798 VDD.t2152 102.87
R6618 VDD.n800 VDD.t1940 102.87
R6619 VDD.n802 VDD.t1878 102.87
R6620 VDD.n809 VDD.t1244 102.87
R6621 VDD.n758 VDD.t1475 102.87
R6622 VDD.n756 VDD.t1679 102.87
R6623 VDD.n834 VDD.t49 102.87
R6624 VDD.n836 VDD.t1081 102.87
R6625 VDD.n838 VDD.t1008 102.87
R6626 VDD.n840 VDD.t1017 102.87
R6627 VDD.n842 VDD.t712 102.87
R6628 VDD.n848 VDD.t1521 102.87
R6629 VDD.n850 VDD.t1558 102.87
R6630 VDD.n852 VDD.t1707 102.87
R6631 VDD.n854 VDD.t1013 102.87
R6632 VDD.n856 VDD.t21 102.87
R6633 VDD.n858 VDD.t1049 102.87
R6634 VDD.n860 VDD.t1944 102.87
R6635 VDD.n866 VDD.t918 102.87
R6636 VDD.n868 VDD.t35 102.87
R6637 VDD.n870 VDD.t1258 102.87
R6638 VDD.n872 VDD.t504 102.87
R6639 VDD.n874 VDD.t710 102.87
R6640 VDD.n881 VDD.t994 102.87
R6641 VDD.n830 VDD.t1356 102.87
R6642 VDD.n828 VDD.t1685 102.87
R6643 VDD.n906 VDD.t650 102.87
R6644 VDD.n908 VDD.t1497 102.87
R6645 VDD.n910 VDD.t783 102.87
R6646 VDD.n912 VDD.t2136 102.87
R6647 VDD.n914 VDD.t618 102.87
R6648 VDD.n920 VDD.t808 102.87
R6649 VDD.n922 VDD.t1626 102.87
R6650 VDD.n924 VDD.t381 102.87
R6651 VDD.n926 VDD.t1283 102.87
R6652 VDD.n928 VDD.t1912 102.87
R6653 VDD.n930 VDD.t670 102.87
R6654 VDD.n932 VDD.t1310 102.87
R6655 VDD.n938 VDD.t749 102.87
R6656 VDD.n940 VDD.t1843 102.87
R6657 VDD.n942 VDD.t1330 102.87
R6658 VDD.n944 VDD.t982 102.87
R6659 VDD.n946 VDD.t2247 102.87
R6660 VDD.n953 VDD.t668 102.87
R6661 VDD.n902 VDD.t532 102.87
R6662 VDD.n900 VDD.t1638 102.87
R6663 VDD.n978 VDD.t771 102.87
R6664 VDD.n980 VDD.t1736 102.87
R6665 VDD.n982 VDD.t39 102.87
R6666 VDD.n984 VDD.t787 102.87
R6667 VDD.n986 VDD.t2100 102.87
R6668 VDD.n992 VDD.t761 102.87
R6669 VDD.n994 VDD.t800 102.87
R6670 VDD.n996 VDD.t393 102.87
R6671 VDD.n998 VDD.t806 102.87
R6672 VDD.n1000 VDD.t1859 102.87
R6673 VDD.n1002 VDD.t759 102.87
R6674 VDD.n1004 VDD.t27 102.87
R6675 VDD.n1010 VDD.t2102 102.87
R6676 VDD.n1012 VDD.t1493 102.87
R6677 VDD.n1014 VDD.t966 102.87
R6678 VDD.n1016 VDD.t1585 102.87
R6679 VDD.n1018 VDD.t580 102.87
R6680 VDD.n1025 VDD.t1035 102.87
R6681 VDD.n974 VDD.t1722 102.87
R6682 VDD.n972 VDD.t444 102.87
R6683 VDD.n1050 VDD.t2162 102.87
R6684 VDD.n1052 VDD.t912 102.87
R6685 VDD.n1054 VDD.t436 102.87
R6686 VDD.n1056 VDD.t1300 102.87
R6687 VDD.n1058 VDD.t1362 102.87
R6688 VDD.n1064 VDD.t2172 102.87
R6689 VDD.n1066 VDD.t1954 102.87
R6690 VDD.n1068 VDD.t67 102.87
R6691 VDD.n1070 VDD.t15 102.87
R6692 VDD.n1072 VDD.t1714 102.87
R6693 VDD.n1074 VDD.t2170 102.87
R6694 VDD.n1076 VDD.t482 102.87
R6695 VDD.n1082 VDD.t1754 102.87
R6696 VDD.n1084 VDD.t940 102.87
R6697 VDD.n1086 VDD.t408 102.87
R6698 VDD.n1088 VDD.t448 102.87
R6699 VDD.n1090 VDD.t1687 102.87
R6700 VDD.n1097 VDD.t2108 102.87
R6701 VDD.n1046 VDD.t71 102.87
R6702 VDD.n1044 VDD.t2178 102.87
R6703 VDD.n1122 VDD.t684 102.87
R6704 VDD.n1124 VDD.t606 102.87
R6705 VDD.n1126 VDD.t1534 102.87
R6706 VDD.n1128 VDD.t952 102.87
R6707 VDD.n1130 VDD.t2116 102.87
R6708 VDD.n1136 VDD.t41 102.87
R6709 VDD.n1138 VDD.t590 102.87
R6710 VDD.n1140 VDD.t2150 102.87
R6711 VDD.n1142 VDD.t486 102.87
R6712 VDD.n1144 VDD.t508 102.87
R6713 VDD.n1146 VDD.t1250 102.87
R6714 VDD.n1148 VDD.t854 102.87
R6715 VDD.n1154 VDD.t960 102.87
R6716 VDD.n1156 VDD.t1542 102.87
R6717 VDD.n1158 VDD.t1279 102.87
R6718 VDD.n1160 VDD.t838 102.87
R6719 VDD.n1162 VDD.t1573 102.87
R6720 VDD.n1169 VDD.t1607 102.87
R6721 VDD.n1118 VDD.t1930 102.87
R6722 VDD.n1116 VDD.t2219 102.87
R6723 VDD.n1194 VDD.t1015 102.87
R6724 VDD.n1196 VDD.t1962 102.87
R6725 VDD.n1198 VDD.t818 102.87
R6726 VDD.n1200 VDD.t1103 102.87
R6727 VDD.n1202 VDD.t47 102.87
R6728 VDD.n1208 VDD.t1473 102.87
R6729 VDD.n1210 VDD.t1886 102.87
R6730 VDD.n1212 VDD.t1896 102.87
R6731 VDD.n1214 VDD.t1304 102.87
R6732 VDD.n1216 VDD.t622 102.87
R6733 VDD.n1218 VDD.t562 102.87
R6734 VDD.n1220 VDD.t954 102.87
R6735 VDD.n1226 VDD.t890 102.87
R6736 VDD.n1228 VDD.t2265 102.87
R6737 VDD.n1230 VDD.t816 102.87
R6738 VDD.n1232 VDD.t2211 102.87
R6739 VDD.n1234 VDD.t690 102.87
R6740 VDD.n1241 VDD.t584 102.87
R6741 VDD.n1190 VDD.t1986 102.87
R6742 VDD.n1188 VDD.t2215 102.87
R6743 VDD.n1266 VDD.t996 102.87
R6744 VDD.n1268 VDD.t1734 102.87
R6745 VDD.n1270 VDD.t656 102.87
R6746 VDD.n1272 VDD.t1804 102.87
R6747 VDD.n1274 VDD.t458 102.87
R6748 VDD.n1280 VDD.t1709 102.87
R6749 VDD.n1282 VDD.t1796 102.87
R6750 VDD.n1284 VDD.t1540 102.87
R6751 VDD.n1286 VDD.t383 102.87
R6752 VDD.n1288 VDD.t51 102.87
R6753 VDD.n1290 VDD.t1603 102.87
R6754 VDD.n1292 VDD.t1471 102.87
R6755 VDD.n1298 VDD.t355 102.87
R6756 VDD.n1300 VDD.t1287 102.87
R6757 VDD.n1302 VDD.t2148 102.87
R6758 VDD.n1304 VDD.t2269 102.87
R6759 VDD.n1306 VDD.t414 102.87
R6760 VDD.n1313 VDD.t1845 102.87
R6761 VDD.n1262 VDD.t602 102.87
R6762 VDD.n1260 VDD.t1926 102.87
R6763 VDD.n1338 VDD.t826 102.87
R6764 VDD.n1340 VDD.t43 102.87
R6765 VDD.n1342 VDD.t1938 102.87
R6766 VDD.n1344 VDD.t1738 102.87
R6767 VDD.n1346 VDD.t2253 102.87
R6768 VDD.n1352 VDD.t654 102.87
R6769 VDD.n1354 VDD.t1732 102.87
R6770 VDD.n1356 VDD.t1861 102.87
R6771 VDD.n1358 VDD.t1589 102.87
R6772 VDD.n1360 VDD.t1616 102.87
R6773 VDD.n1362 VDD.t578 102.87
R6774 VDD.n1364 VDD.t1587 102.87
R6775 VDD.n1370 VDD.t1770 102.87
R6776 VDD.n1372 VDD.t81 102.87
R6777 VDD.n1374 VDD.t2094 102.87
R6778 VDD.n1376 VDD.t1664 102.87
R6779 VDD.n1378 VDD.t1265 102.87
R6780 VDD.n1385 VDD.t1517 102.87
R6781 VDD.n1334 VDD.t984 102.87
R6782 VDD.n1332 VDD.t2144 102.87
R6783 VDD.n1410 VDD.t1898 102.87
R6784 VDD.n1412 VDD.t1000 102.87
R6785 VDD.n1414 VDD.t886 102.87
R6786 VDD.n1416 VDD.t476 102.87
R6787 VDD.n1418 VDD.t1652 102.87
R6788 VDD.n1424 VDD.t468 102.87
R6789 VDD.n1426 VDD.t600 102.87
R6790 VDD.n1428 VDD.t2234 102.87
R6791 VDD.n1430 VDD.t1461 102.87
R6792 VDD.n1432 VDD.t914 102.87
R6793 VDD.n1434 VDD.t1705 102.87
R6794 VDD.n1436 VDD.t341 102.87
R6795 VDD.n1442 VDD.t2002 102.87
R6796 VDD.n1444 VDD.t990 102.87
R6797 VDD.n1446 VDD.t1546 102.87
R6798 VDD.n1448 VDD.t1874 102.87
R6799 VDD.n1450 VDD.t311 102.87
R6800 VDD.n1457 VDD.t1564 102.87
R6801 VDD.n1406 VDD.t948 102.87
R6802 VDD.n1404 VDD.t540 102.87
R6803 VDD.n1482 VDD.t1847 102.87
R6804 VDD.n1484 VDD.t1099 102.87
R6805 VDD.n1486 VDD.t1666 102.87
R6806 VDD.n1488 VDD.t331 102.87
R6807 VDD.n1490 VDD.t359 102.87
R6808 VDD.n1496 VDD.t1281 102.87
R6809 VDD.n1498 VDD.t832 102.87
R6810 VDD.n1500 VDD.t946 102.87
R6811 VDD.n1502 VDD.t1560 102.87
R6812 VDD.n1504 VDD.t1386 102.87
R6813 VDD.n1506 VDD.t1849 102.87
R6814 VDD.n1508 VDD.t1409 102.87
R6815 VDD.n1514 VDD.t1746 102.87
R6816 VDD.n1516 VDD.t1837 102.87
R6817 VDD.n1518 VDD.t904 102.87
R6818 VDD.n1520 VDD.t1865 102.87
R6819 VDD.n1522 VDD.t1599 102.87
R6820 VDD.n1529 VDD.t450 102.87
R6821 VDD.n1478 VDD.t524 102.87
R6822 VDD.n1476 VDD.t2130 102.87
R6823 VDD.n1554 VDD.t1324 102.87
R6824 VDD.n1556 VDD.t1469 102.87
R6825 VDD.n1558 VDD.t930 102.87
R6826 VDD.n1560 VDD.t2209 102.87
R6827 VDD.n1562 VDD.t2236 102.87
R6828 VDD.n1568 VDD.t1232 102.87
R6829 VDD.n1570 VDD.t1827 102.87
R6830 VDD.n1572 VDD.t1340 102.87
R6831 VDD.n1574 VDD.t379 102.87
R6832 VDD.n1576 VDD.t658 102.87
R6833 VDD.n1578 VDD.t2112 102.87
R6834 VDD.n1580 VDD.t755 102.87
R6835 VDD.n1586 VDD.t588 102.87
R6836 VDD.n1588 VDD.t598 102.87
R6837 VDD.n1590 VDD.t1025 102.87
R6838 VDD.n1592 VDD.t534 102.87
R6839 VDD.n1594 VDD.t1752 102.87
R6840 VDD.n1601 VDD.t810 102.87
R6841 VDD.n1550 VDD.t1634 102.87
R6842 VDD.n1548 VDD.t1726 102.87
R6843 VDD.n1674 VDD.t1275 102.87
R6844 VDD.n1670 VDD.t958 102.87
R6845 VDD.n1668 VDD.t1992 102.87
R6846 VDD.n1666 VDD.t1946 102.87
R6847 VDD.n1664 VDD.t1900 102.87
R6848 VDD.n1662 VDD.t644 102.87
R6849 VDD.n1658 VDD.t353 102.87
R6850 VDD.n1656 VDD.t680 102.87
R6851 VDD.n1654 VDD.t418 102.87
R6852 VDD.n1652 VDD.t396 102.87
R6853 VDD.n1650 VDD.t1876 102.87
R6854 VDD.n1648 VDD.t564 102.87
R6855 VDD.n1646 VDD.t323 102.87
R6856 VDD.n1642 VDD.t1994 102.87
R6857 VDD.n1640 VDD.t387 102.87
R6858 VDD.n1638 VDD.t1672 102.87
R6859 VDD.n1636 VDD.t678 102.87
R6860 VDD.n1634 VDD.t2281 102.87
R6861 VDD.n1630 VDD.t696 102.87
R6862 VDD.n1628 VDD.t822 102.87
R6863 VDD.n586 VDD.t1033 102.87
R6864 VDD.n584 VDD.t928 102.87
R6865 VDD.n582 VDD.t840 102.87
R6866 VDD.n580 VDD.t1065 102.87
R6867 VDD.n578 VDD.t864 102.87
R6868 VDD.n574 VDD.t1918 102.87
R6869 VDD.n572 VDD.t1051 102.87
R6870 VDD.n570 VDD.t1618 102.87
R6871 VDD.n568 VDD.t357 102.87
R6872 VDD.n566 VDD.t347 102.87
R6873 VDD.n564 VDD.t1910 102.87
R6874 VDD.n562 VDD.t478 102.87
R6875 VDD.n558 VDD.t740 102.87
R6876 VDD.n556 VDD.t373 102.87
R6877 VDD.n554 VDD.t1390 102.87
R6878 VDD.n552 VDD.t2232 102.87
R6879 VDD.n550 VDD.t1774 102.87
R6880 VDD.n546 VDD.t2124 102.87
R6881 VDD.n544 VDD.t2229 102.87
R6882 VDD.n609 VDD.t698 102.87
R6883 VDD.n611 VDD.t1175 102.87
R6884 VDD.n618 VDD.t936 102.87
R6885 VDD.n620 VDD.t75 102.87
R6886 VDD.n622 VDD.t1683 102.87
R6887 VDD.n624 VDD.t574 102.87
R6888 VDD.n626 VDD.t538 102.87
R6889 VDD.n632 VDD.t1872 102.87
R6890 VDD.n634 VDD.t732 102.87
R6891 VDD.n636 VDD.t660 102.87
R6892 VDD.n638 VDD.t1964 102.87
R6893 VDD.n640 VDD.t718 102.87
R6894 VDD.n642 VDD.t888 102.87
R6895 VDD.n644 VDD.t1695 102.87
R6896 VDD.n650 VDD.t333 102.87
R6897 VDD.n652 VDD.t1047 102.87
R6898 VDD.n654 VDD.t910 102.87
R6899 VDD.n656 VDD.t1093 102.87
R6900 VDD.n658 VDD.t852 102.87
R6901 VDD.n665 VDD.t1503 102.87
R6902 VDD.n593 VDD.t2285 102.87
R6903 VDD.n701 VDD.t2255 98.665
R6904 VDD.n719 VDD.t1609 98.665
R6905 VDD.n672 VDD.t1487 98.665
R6906 VDD.n773 VDD.t1792 98.665
R6907 VDD.n791 VDD.t765 98.665
R6908 VDD.n744 VDD.t1906 98.665
R6909 VDD.n845 VDD.t1 98.665
R6910 VDD.n863 VDD.t1191 98.665
R6911 VDD.n816 VDD.t2273 98.665
R6912 VDD.n917 VDD.t2004 98.665
R6913 VDD.n935 VDD.t484 98.665
R6914 VDD.n888 VDD.t1670 98.665
R6915 VDD.n989 VDD.t1077 98.665
R6916 VDD.n1007 VDD.t2118 98.665
R6917 VDD.n960 VDD.t1888 98.665
R6918 VDD.n1061 VDD.t1811 98.665
R6919 VDD.n1079 VDD.t576 98.665
R6920 VDD.n1032 VDD.t1740 98.665
R6921 VDD.n1133 VDD.t1863 98.665
R6922 VDD.n1151 VDD.t868 98.665
R6923 VDD.n1104 VDD.t1346 98.665
R6924 VDD.n1205 VDD.t11 98.665
R6925 VDD.n1223 VDD.t1374 98.665
R6926 VDD.n1176 VDD.t2182 98.665
R6927 VDD.n1277 VDD.t926 98.665
R6928 VDD.n1295 VDD.t1570 98.665
R6929 VDD.n1248 VDD.t315 98.665
R6930 VDD.n1349 VDD.t1650 98.665
R6931 VDD.n1367 VDD.t1972 98.665
R6932 VDD.n1320 VDD.t1934 98.665
R6933 VDD.n1421 VDD.t526 98.665
R6934 VDD.n1439 VDD.t1784 98.665
R6935 VDD.n1392 VDD.t1756 98.665
R6936 VDD.n1493 VDD.t612 98.665
R6937 VDD.n1511 VDD.t1234 98.665
R6938 VDD.n1464 VDD.t3 98.665
R6939 VDD.n1565 VDD.t500 98.665
R6940 VDD.n1583 VDD.t922 98.665
R6941 VDD.n1536 VDD.t1402 98.665
R6942 VDD.n1609 VDD.t1984 98.665
R6943 VDD.n1611 VDD.t446 98.665
R6944 VDD.n1613 VDD.t844 98.665
R6945 VDD.n1616 VDD.t2000 98.665
R6946 VDD.n528 VDD.t1302 98.665
R6947 VDD.n530 VDD.t422 98.665
R6948 VDD.n533 VDD.t1432 98.665
R6949 VDD.n615 VDD.t1902 98.665
R6950 VDD.n629 VDD.t1924 98.665
R6951 VDD.n647 VDD.t1855 98.665
R6952 VDD.n590 VDD.t1067 98.665
R6953 VDD.n734 VDD.t1087 98.665
R6954 VDD.n806 VDD.t1622 98.665
R6955 VDD.n878 VDD.t722 98.665
R6956 VDD.n950 VDD.t964 98.665
R6957 VDD.n1022 VDD.t542 98.665
R6958 VDD.n1094 VDD.t57 98.665
R6959 VDD.n1166 VDD.t2197 98.665
R6960 VDD.n1238 VDD.t676 98.665
R6961 VDD.n1310 VDD.t1817 98.665
R6962 VDD.n1382 VDD.t1436 98.665
R6963 VDD.n1454 VDD.t708 98.665
R6964 VDD.n1526 VDD.t751 98.665
R6965 VDD.n1598 VDD.t2193 98.665
R6966 VDD.n662 VDD.t1642 98.665
R6967 VDD.t364 VDD.t362 96.694
R6968 VDD.t425 VDD.t1044 96.694
R6969 VDD.t1775 VDD.t1590 96.694
R6970 VDD.t827 VDD.t1270 96.694
R6971 VDD.t746 VDD.t797 96.694
R6972 VDD.t1054 VDD.t401 96.694
R6973 VDD.t1227 VDD.t1084 96.694
R6974 VDD.t471 VDD.t979 96.694
R6975 VDD.t1673 VDD.t623 96.694
R6976 VDD.t22 VDD.t72 96.694
R6977 VDD.t1429 VDD.t1655 96.694
R6978 VDD.t1276 VDD.t1508 96.694
R6979 VDD.t32 VDD.t60 96.694
R6980 VDD.t1237 VDD.t565 96.694
R6981 VDD.t18 VDD.t1036 96.694
R6982 VDD.t681 VDD.t877 95.697
R6983 VDD.n680 VDD.t1220 86.102
R6984 VDD.n824 VDD.t1198 86.102
R6985 VDD.n968 VDD.t1194 86.102
R6986 VDD.n1112 VDD.t1206 86.102
R6987 VDD.n1256 VDD.t1202 86.102
R6988 VDD.n1400 VDD.t1218 86.102
R6989 VDD.n540 VDD.t1212 86.102
R6990 VDD.n1544 VDD.t1216 86.057
R6991 VDD.n118 VDD.t114 85.729
R6992 VDD.n150 VDD.t194 85.729
R6993 VDD.n182 VDD.t198 85.729
R6994 VDD.n214 VDD.t118 85.729
R6995 VDD.n246 VDD.t138 85.729
R6996 VDD.n278 VDD.t176 85.729
R6997 VDD.n310 VDD.t120 85.729
R6998 VDD.n342 VDD.t128 85.729
R6999 VDD.n374 VDD.t146 85.729
R7000 VDD.n406 VDD.t214 85.729
R7001 VDD.n438 VDD.t168 85.729
R7002 VDD.n470 VDD.t158 85.729
R7003 VDD.n502 VDD.t92 85.729
R7004 VDD.n752 VDD.t1214 85.525
R7005 VDD.n896 VDD.t1210 85.525
R7006 VDD.n1040 VDD.t1224 85.525
R7007 VDD.n1184 VDD.t1196 85.525
R7008 VDD.n1328 VDD.t1208 85.525
R7009 VDD.n1472 VDD.t1204 85.525
R7010 VDD.n605 VDD.t1200 85.525
R7011 VDD.n689 VDD.t1701 85.516
R7012 VDD.n691 VDD.t1970 85.516
R7013 VDD.n693 VDD.t1758 85.516
R7014 VDD.n695 VDD.t972 85.516
R7015 VDD.n697 VDD.t548 85.516
R7016 VDD.n699 VDD.t986 85.516
R7017 VDD.n703 VDD.t2283 85.516
R7018 VDD.n705 VDD.t462 85.516
R7019 VDD.n707 VDD.t2008 85.516
R7020 VDD.n709 VDD.t769 85.516
R7021 VDD.n711 VDD.t842 85.516
R7022 VDD.n713 VDD.t1748 85.516
R7023 VDD.n715 VDD.t536 85.516
R7024 VDD.n717 VDD.t1548 85.516
R7025 VDD.n721 VDD.t880 85.516
R7026 VDD.n723 VDD.t339 85.516
R7027 VDD.n725 VDD.t2126 85.516
R7028 VDD.n727 VDD.t1605 85.516
R7029 VDD.n729 VDD.t2164 85.516
R7030 VDD.n731 VDD.t898 85.516
R7031 VDD.n738 VDD.t1411 85.516
R7032 VDD.n736 VDD.t944 85.516
R7033 VDD.n687 VDD.t1841 85.516
R7034 VDD.n685 VDD.t2203 85.516
R7035 VDD.n761 VDD.t1974 85.516
R7036 VDD.n763 VDD.t2158 85.516
R7037 VDD.n765 VDD.t634 85.516
R7038 VDD.n767 VDD.t59 85.516
R7039 VDD.n769 VDD.t1942 85.516
R7040 VDD.n771 VDD.t1428 85.516
R7041 VDD.n775 VDD.t1636 85.516
R7042 VDD.n777 VDD.t1171 85.516
R7043 VDD.n779 VDD.t440 85.516
R7044 VDD.n781 VDD.t777 85.516
R7045 VDD.n783 VDD.t1800 85.516
R7046 VDD.n785 VDD.t2238 85.516
R7047 VDD.n787 VDD.t2180 85.516
R7048 VDD.n789 VDD.t351 85.516
R7049 VDD.n793 VDD.t1483 85.516
R7050 VDD.n795 VDD.t522 85.516
R7051 VDD.n797 VDD.t412 85.516
R7052 VDD.n799 VDD.t2146 85.516
R7053 VDD.n801 VDD.t2006 85.516
R7054 VDD.n803 VDD.t1880 85.516
R7055 VDD.n810 VDD.t570 85.516
R7056 VDD.n808 VDD.t385 85.516
R7057 VDD.n759 VDD.t1479 85.516
R7058 VDD.n757 VDD.t1459 85.516
R7059 VDD.n833 VDD.t2275 85.516
R7060 VDD.n835 VDD.t45 85.516
R7061 VDD.n837 VDD.t1079 85.516
R7062 VDD.n839 VDD.t369 85.516
R7063 VDD.n841 VDD.t2132 85.516
R7064 VDD.n843 VDD.t702 85.516
R7065 VDD.n847 VDD.t1691 85.516
R7066 VDD.n849 VDD.t652 85.516
R7067 VDD.n851 VDD.t1632 85.516
R7068 VDD.n853 VDD.t694 85.516
R7069 VDD.n855 VDD.t1562 85.516
R7070 VDD.n857 VDD.t9 85.516
R7071 VDD.n859 VDD.t434 85.516
R7072 VDD.n861 VDD.t2120 85.516
R7073 VDD.n865 VDD.t610 85.516
R7074 VDD.n867 VDD.t1312 85.516
R7075 VDD.n869 VDD.t25 85.516
R7076 VDD.n871 VDD.t1703 85.516
R7077 VDD.n873 VDD.t2140 85.516
R7078 VDD.n875 VDD.t1904 85.516
R7079 VDD.n882 VDD.t866 85.516
R7080 VDD.n880 VDD.t1465 85.516
R7081 VDD.n831 VDD.t1358 85.516
R7082 VDD.n829 VDD.t830 85.516
R7083 VDD.n905 VDD.t1658 85.516
R7084 VDD.n907 VDD.t648 85.516
R7085 VDD.n909 VDD.t1463 85.516
R7086 VDD.n911 VDD.t892 85.516
R7087 VDD.n913 VDD.t2249 85.516
R7088 VDD.n915 VDD.t640 85.516
R7089 VDD.n919 VDD.t1988 85.516
R7090 VDD.n921 VDD.t796 85.516
R7091 VDD.n923 VDD.t608 85.516
R7092 VDD.n925 VDD.t530 85.516
R7093 VDD.n927 VDD.t1813 85.516
R7094 VDD.n929 VDD.t1720 85.516
R7095 VDD.n931 VDD.t1230 85.516
R7096 VDD.n933 VDD.t1491 85.516
R7097 VDD.n937 VDD.t1697 85.516
R7098 VDD.n939 VDD.t1248 85.516
R7099 VDD.n941 VDD.t773 85.516
R7100 VDD.n943 VDD.t1819 85.516
R7101 VDD.n945 VDD.t456 85.516
R7102 VDD.n947 VDD.t2227 85.516
R7103 VDD.n954 VDD.t1867 85.516
R7104 VDD.n952 VDD.t962 85.516
R7105 VDD.n903 VDD.t1326 85.516
R7106 VDD.n901 VDD.t1624 85.516
R7107 VDD.n977 VDD.t779 85.516
R7108 VDD.n979 VDD.t726 85.516
R7109 VDD.n981 VDD.t1515 85.516
R7110 VDD.n983 VDD.t53 85.516
R7111 VDD.n985 VDD.t1831 85.516
R7112 VDD.n987 VDD.t2251 85.516
R7113 VDD.n991 VDD.t460 85.516
R7114 VDD.n993 VDD.t1328 85.516
R7115 VDD.n995 VDD.t1566 85.516
R7116 VDD.n997 VDD.t430 85.516
R7117 VDD.n999 VDD.t1424 85.516
R7118 VDD.n1001 VDD.t970 85.516
R7119 VDD.n1003 VDD.t1839 85.516
R7120 VDD.n1005 VDD.t745 85.516
R7121 VDD.n1009 VDD.t932 85.516
R7122 VDD.n1011 VDD.t410 85.516
R7123 VDD.n1013 VDD.t672 85.516
R7124 VDD.n1015 VDD.t1398 85.516
R7125 VDD.n1017 VDD.t1370 85.516
R7126 VDD.n1019 VDD.t582 85.516
R7127 VDD.n1026 VDD.t345 85.516
R7128 VDD.n1024 VDD.t1344 85.516
R7129 VDD.n975 VDD.t1376 85.516
R7130 VDD.n973 VDD.t1760 85.516
R7131 VDD.n1049 VDD.t730 85.516
R7132 VDD.n1051 VDD.t616 85.516
R7133 VDD.n1053 VDD.t1246 85.516
R7134 VDD.n1055 VDD.t1360 85.516
R7135 VDD.n1057 VDD.t1298 85.516
R7136 VDD.n1059 VDD.t1364 85.516
R7137 VDD.n1063 VDD.t1762 85.516
R7138 VDD.n1065 VDD.t13 85.516
R7139 VDD.n1067 VDD.t1960 85.516
R7140 VDD.n1069 VDD.t83 85.516
R7141 VDD.n1071 VDD.t1544 85.516
R7142 VDD.n1073 VDD.t1716 85.516
R7143 VDD.n1075 VDD.t1267 85.516
R7144 VDD.n1077 VDD.t452 85.516
R7145 VDD.n1081 VDD.t560 85.516
R7146 VDD.n1083 VDD.t377 85.516
R7147 VDD.n1085 VDD.t942 85.516
R7148 VDD.n1087 VDD.t391 85.516
R7149 VDD.n1089 VDD.t1495 85.516
R7150 VDD.n1091 VDD.t1718 85.516
R7151 VDD.n1098 VDD.t2257 85.516
R7152 VDD.n1096 VDD.t2201 85.516
R7153 VDD.n1047 VDD.t37 85.516
R7154 VDD.n1045 VDD.t2185 85.516
R7155 VDD.n1121 VDD.t662 85.516
R7156 VDD.n1123 VDD.t1314 85.516
R7157 VDD.n1125 VDD.t1256 85.516
R7158 VDD.n1127 VDD.t1029 85.516
R7159 VDD.n1129 VDD.t1378 85.516
R7160 VDD.n1131 VDD.t2104 85.516
R7161 VDD.n1135 VDD.t2122 85.516
R7162 VDD.n1137 VDD.t2189 85.516
R7163 VDD.n1139 VDD.t1595 85.516
R7164 VDD.n1141 VDD.t321 85.516
R7165 VDD.n1143 VDD.t1612 85.516
R7166 VDD.n1145 VDD.t466 85.516
R7167 VDD.n1147 VDD.t908 85.516
R7168 VDD.n1149 VDD.t1786 85.516
R7169 VDD.n1153 VDD.t992 85.516
R7170 VDD.n1155 VDD.t1681 85.516
R7171 VDD.n1157 VDD.t1260 85.516
R7172 VDD.n1159 VDD.t1332 85.516
R7173 VDD.n1161 VDD.t1189 85.516
R7174 VDD.n1163 VDD.t1870 85.516
R7175 VDD.n1170 VDD.t988 85.516
R7176 VDD.n1168 VDD.t2207 85.516
R7177 VDD.n1119 VDD.t55 85.516
R7178 VDD.n1117 VDD.t2213 85.516
R7179 VDD.n1193 VDD.t2168 85.516
R7180 VDD.n1195 VDD.t1426 85.516
R7181 VDD.n1197 VDD.t1956 85.516
R7182 VDD.n1199 VDD.t792 85.516
R7183 VDD.n1201 VDD.t1101 85.516
R7184 VDD.n1203 VDD.t85 85.516
R7185 VDD.n1207 VDD.t7 85.516
R7186 VDD.n1209 VDD.t1477 85.516
R7187 VDD.n1211 VDD.t520 85.516
R7188 VDD.n1213 VDD.t950 85.516
R7189 VDD.n1215 VDD.t1392 85.516
R7190 VDD.n1217 VDD.t361 85.516
R7191 VDD.n1219 VDD.t517 85.516
R7192 VDD.n1221 VDD.t688 85.516
R7193 VDD.n1225 VDD.t1772 85.516
R7194 VDD.n1227 VDD.t1768 85.516
R7195 VDD.n1229 VDD.t2267 85.516
R7196 VDD.n1231 VDD.t2187 85.516
R7197 VDD.n1233 VDD.t2221 85.516
R7198 VDD.n1235 VDD.t686 85.516
R7199 VDD.n1242 VDD.t1027 85.516
R7200 VDD.n1240 VDD.t674 85.516
R7201 VDD.n1191 VDD.t1920 85.516
R7202 VDD.n1189 VDD.t2199 85.516
R7203 VDD.n1265 VDD.t313 85.516
R7204 VDD.n1267 VDD.t2223 85.516
R7205 VDD.n1269 VDD.t1806 85.516
R7206 VDD.n1271 VDD.t586 85.516
R7207 VDD.n1273 VDD.t1802 85.516
R7208 VDD.n1275 VDD.t1352 85.516
R7209 VDD.n1279 VDD.t1368 85.516
R7210 VDD.n1281 VDD.t424 85.516
R7211 VDD.n1283 VDD.t1821 85.516
R7212 VDD.n1285 VDD.t596 85.516
R7213 VDD.n1287 VDD.t956 85.516
R7214 VDD.n1289 VDD.t319 85.516
R7215 VDD.n1291 VDD.t1614 85.516
R7216 VDD.n1293 VDD.t1057 85.516
R7217 VDD.n1297 VDD.t628 85.516
R7218 VDD.n1299 VDD.t1575 85.516
R7219 VDD.n1301 VDD.t2217 85.516
R7220 VDD.n1303 VDD.t329 85.516
R7221 VDD.n1305 VDD.t2174 85.516
R7222 VDD.n1307 VDD.t506 85.516
R7223 VDD.n1314 VDD.t464 85.516
R7224 VDD.n1312 VDD.t1481 85.516
R7225 VDD.n1263 VDD.t604 85.516
R7226 VDD.n1261 VDD.t1922 85.516
R7227 VDD.n1337 VDD.t2154 85.516
R7228 VDD.n1339 VDD.t814 85.516
R7229 VDD.n1341 VDD.t65 85.516
R7230 VDD.n1343 VDD.t1936 85.516
R7231 VDD.n1345 VDD.t442 85.516
R7232 VDD.n1347 VDD.t757 85.516
R7233 VDD.n1351 VDD.t1648 85.516
R7234 VDD.n1353 VDD.t528 85.516
R7235 VDD.n1355 VDD.t371 85.516
R7236 VDD.n1357 VDD.t642 85.516
R7237 VDD.n1359 VDD.t1059 85.516
R7238 VDD.n1361 VDD.t1829 85.516
R7239 VDD.n1363 VDD.t550 85.516
R7240 VDD.n1365 VDD.t568 85.516
R7241 VDD.n1369 VDD.t1908 85.516
R7242 VDD.n1371 VDD.t1778 85.516
R7243 VDD.n1373 VDD.t1660 85.516
R7244 VDD.n1375 VDD.t1968 85.516
R7245 VDD.n1377 VDD.t1662 85.516
R7246 VDD.n1379 VDD.t692 85.516
R7247 VDD.n1386 VDD.t1523 85.516
R7248 VDD.n1384 VDD.t594 85.516
R7249 VDD.n1335 VDD.t1396 85.516
R7250 VDD.n1333 VDD.t1914 85.516
R7251 VDD.n1409 VDD.t1348 85.516
R7252 VDD.n1411 VDD.t1894 85.516
R7253 VDD.n1413 VDD.t1002 85.516
R7254 VDD.n1415 VDD.t1780 85.516
R7255 VDD.n1417 VDD.t1226 85.516
R7256 VDD.n1419 VDD.t592 85.516
R7257 VDD.n1423 VDD.t1527 85.516
R7258 VDD.n1425 VDD.t389 85.516
R7259 VDD.n1427 VDD.t1418 85.516
R7260 VDD.n1429 VDD.t2242 85.516
R7261 VDD.n1431 VDD.t1794 85.516
R7262 VDD.n1433 VDD.t1513 85.516
R7263 VDD.n1435 VDD.t876 85.516
R7264 VDD.n1437 VDD.t1262 85.516
R7265 VDD.n1441 VDD.t858 85.516
R7266 VDD.n1443 VDD.t1990 85.516
R7267 VDD.n1445 VDD.t488 85.516
R7268 VDD.n1447 VDD.t1742 85.516
R7269 VDD.n1449 VDD.t870 85.516
R7270 VDD.n1451 VDD.t317 85.516
R7271 VDD.n1458 VDD.t496 85.516
R7272 VDD.n1456 VDD.t1269 85.516
R7273 VDD.n1407 VDD.t400 85.516
R7274 VDD.n1405 VDD.t1011 85.516
R7275 VDD.n1481 VDD.t1519 85.516
R7276 VDD.n1483 VDD.t1525 85.516
R7277 VDD.n1485 VDD.t734 85.516
R7278 VDD.n1487 VDD.t924 85.516
R7279 VDD.n1489 VDD.t1285 85.516
R7280 VDD.n1491 VDD.t934 85.516
R7281 VDD.n1495 VDD.t706 85.516
R7282 VDD.n1497 VDD.t1306 85.516
R7283 VDD.n1499 VDD.t834 85.516
R7284 VDD.n1501 VDD.t1579 85.516
R7285 VDD.n1503 VDD.t494 85.516
R7286 VDD.n1505 VDD.t1384 85.516
R7287 VDD.n1507 VDD.t1422 85.516
R7288 VDD.n1509 VDD.t1407 85.516
R7289 VDD.n1513 VDD.t546 85.516
R7290 VDD.n1515 VDD.t1489 85.516
R7291 VDD.n1517 VDD.t1689 85.516
R7292 VDD.n1519 VDD.t1091 85.516
R7293 VDD.n1521 VDD.t1744 85.516
R7294 VDD.n1523 VDD.t1043 85.516
R7295 VDD.n1530 VDD.t1380 85.516
R7296 VDD.n1528 VDD.t1273 85.516
R7297 VDD.n1479 VDD.t1179 85.516
R7298 VDD.n1477 VDD.t1952 85.516
R7299 VDD.n1553 VDD.t976 85.516
R7300 VDD.n1555 VDD.t1322 85.516
R7301 VDD.n1557 VDD.t1350 85.516
R7302 VDD.n1559 VDD.t1976 85.516
R7303 VDD.n1561 VDD.t2191 85.516
R7304 VDD.n1563 VDD.t882 85.516
R7305 VDD.n1567 VDD.t1293 85.516
R7306 VDD.n1569 VDD.t1628 85.516
R7307 VDD.n1571 VDD.t820 85.516
R7308 VDD.n1573 VDD.t1342 85.516
R7309 VDD.n1575 VDD.t1413 85.516
R7310 VDD.n1577 VDD.t1892 85.516
R7311 VDD.n1579 VDD.t2114 85.516
R7312 VDD.n1581 VDD.t1499 85.516
R7313 VDD.n1585 VDD.t416 85.516
R7314 VDD.n1587 VDD.t1825 85.516
R7315 VDD.n1589 VDD.t1556 85.516
R7316 VDD.n1591 VDD.t1021 85.516
R7317 VDD.n1593 VDD.t515 85.516
R7318 VDD.n1595 VDD.t1187 85.516
R7319 VDD.n1602 VDD.t736 85.516
R7320 VDD.n1600 VDD.t17 85.516
R7321 VDD.n1551 VDD.t1501 85.516
R7322 VDD.n1549 VDD.t1724 85.516
R7323 VDD.n1675 VDD.t632 85.516
R7324 VDD.n1673 VDD.t1928 85.516
R7325 VDD.n1671 VDD.t1577 85.516
R7326 VDD.n1669 VDD.t2134 85.516
R7327 VDD.n1667 VDD.t1950 85.516
R7328 VDD.n1665 VDD.t2098 85.516
R7329 VDD.n1663 VDD.t1438 85.516
R7330 VDD.n1661 VDD.t763 85.516
R7331 VDD.n1659 VDD.t1075 85.516
R7332 VDD.n1657 VDD.t1405 85.516
R7333 VDD.n1655 VDD.t406 85.516
R7334 VDD.n1653 VDD.t404 85.516
R7335 VDD.n1651 VDD.t1240 85.516
R7336 VDD.n1649 VDD.t1440 85.516
R7337 VDD.n1647 VDD.t325 85.516
R7338 VDD.n1645 VDD.t1334 85.516
R7339 VDD.n1643 VDD.t2244 85.516
R7340 VDD.n1641 VDD.t1529 85.516
R7341 VDD.n1639 VDD.t1454 85.516
R7342 VDD.n1637 VDD.t900 85.516
R7343 VDD.n1635 VDD.t2010 85.516
R7344 VDD.n1633 VDD.t2138 85.516
R7345 VDD.n1631 VDD.t558 85.516
R7346 VDD.n1629 VDD.t824 85.516
R7347 VDD.n587 VDD.t1782 85.516
R7348 VDD.n585 VDD.t1630 85.516
R7349 VDD.n583 VDD.t1366 85.516
R7350 VDD.n581 VDD.t704 85.516
R7351 VDD.n579 VDD.t836 85.516
R7352 VDD.n577 VDD.t1039 85.516
R7353 VDD.n575 VDD.t1552 85.516
R7354 VDD.n573 VDD.t502 85.516
R7355 VDD.n571 VDD.t1823 85.516
R7356 VDD.n569 VDD.t480 85.516
R7357 VDD.n567 VDD.t1890 85.516
R7358 VDD.n565 VDD.t2128 85.516
R7359 VDD.n563 VDD.t1809 85.516
R7360 VDD.n561 VDD.t902 85.516
R7361 VDD.n559 VDD.t738 85.516
R7362 VDD.n557 VDD.t375 85.516
R7363 VDD.n555 VDD.t1095 85.516
R7364 VDD.n553 VDD.t2240 85.516
R7365 VDD.n551 VDD.t714 85.516
R7366 VDD.n549 VDD.t1485 85.516
R7367 VDD.n547 VDD.t1948 85.516
R7368 VDD.n545 VDD.t2156 85.516
R7369 VDD.n610 VDD.t1693 85.516
R7370 VDD.n612 VDD.t1958 85.516
R7371 VDD.n617 VDD.t614 85.516
R7372 VDD.n619 VDD.t646 85.516
R7373 VDD.n621 VDD.t69 85.516
R7374 VDD.n623 VDD.t896 85.516
R7375 VDD.n625 VDD.t1583 85.516
R7376 VDD.n627 VDD.t1041 85.516
R7377 VDD.n631 VDD.t1932 85.516
R7378 VDD.n633 VDD.t1996 85.516
R7379 VDD.n635 VDD.t1063 85.516
R7380 VDD.n637 VDD.t1916 85.516
R7381 VDD.n639 VDD.t1730 85.516
R7382 VDD.n641 VDD.t716 85.516
R7383 VDD.n643 VDD.t490 85.516
R7384 VDD.n645 VDD.t906 85.516
R7385 VDD.n649 VDD.t1882 85.516
R7386 VDD.n651 VDD.t79 85.516
R7387 VDD.n653 VDD.t630 85.516
R7388 VDD.n655 VDD.t1415 85.516
R7389 VDD.n657 VDD.t343 85.516
R7390 VDD.n659 VDD.t1668 85.516
R7391 VDD.n666 VDD.t802 85.516
R7392 VDD.n664 VDD.t470 85.516
R7393 VDD.n592 VDD.t856 85.516
R7394 VDD.n594 VDD.t1394 85.516
R7395 VDD.n1624 VDD.t1222 85.47
R7396 VDD.n22 VDD.t106 84.732
R7397 VDD.n54 VDD.t100 84.732
R7398 VDD.n86 VDD.t188 84.732
R7399 VDD.n1678 VDD.n526 73.57
R7400 VDD.n603 VDD.n602 44.423
R7401 VDD.n598 VDD.t1236 34.491
R7402 VDD.n674 VDD.t1790 34.491
R7403 VDD.n746 VDD.t1798 34.491
R7404 VDD.n818 VDD.t572 34.491
R7405 VDD.n890 VDD.t513 34.491
R7406 VDD.n962 VDD.t428 34.491
R7407 VDD.n1034 VDD.t1173 34.491
R7408 VDD.n1106 VDD.t1177 34.491
R7409 VDD.n1178 VDD.t1320 34.491
R7410 VDD.n1250 VDD.t2195 34.491
R7411 VDD.n1322 VDD.t742 34.491
R7412 VDD.n1394 VDD.t327 34.491
R7413 VDD.n1466 VDD.t2259 34.491
R7414 VDD.n1538 VDD.t1699 34.491
R7415 VDD.n1618 VDD.t1183 34.491
R7416 VDD.n535 VDD.t620 34.491
R7417 VDD.n598 VDD.t432 34.259
R7418 VDD.n674 VDD.t1788 34.259
R7419 VDD.n746 VDD.t1982 34.259
R7420 VDD.n818 VDD.t1581 34.259
R7421 VDD.n890 VDD.t31 34.259
R7422 VDD.n962 VDD.t1073 34.259
R7423 VDD.n1034 VDD.t1400 34.259
R7424 VDD.n1106 VDD.t5 34.259
R7425 VDD.n1178 VDD.t1061 34.259
R7426 VDD.n1250 VDD.t337 34.259
R7427 VDD.n1322 VDD.t1457 34.259
R7428 VDD.n1394 VDD.t753 34.259
R7429 VDD.n1466 VDD.t2110 34.259
R7430 VDD.n1538 VDD.t1711 34.259
R7431 VDD.n1618 VDD.t1676 34.259
R7432 VDD.n535 VDD.t1833 34.259
R7433 VDD.n23 VDD.n22 24.245
R7434 VDD.n55 VDD.n54 24.245
R7435 VDD.n87 VDD.n86 24.245
R7436 VDD.n119 VDD.n118 24.245
R7437 VDD.n151 VDD.n150 24.245
R7438 VDD.n183 VDD.n182 24.245
R7439 VDD.n215 VDD.n214 24.245
R7440 VDD.n247 VDD.n246 24.245
R7441 VDD.n279 VDD.n278 24.245
R7442 VDD.n311 VDD.n310 24.245
R7443 VDD.n343 VDD.n342 24.245
R7444 VDD.n375 VDD.n374 24.245
R7445 VDD.n407 VDD.n406 24.245
R7446 VDD.n439 VDD.n438 24.245
R7447 VDD.n471 VDD.n470 24.245
R7448 VDD.n503 VDD.n502 24.245
R7449 VDD.n676 VDD.t1149 20.995
R7450 VDD.n748 VDD.t1157 20.995
R7451 VDD.n820 VDD.t1127 20.995
R7452 VDD.n892 VDD.t1163 20.995
R7453 VDD.n964 VDD.t1119 20.995
R7454 VDD.n1036 VDD.t1139 20.995
R7455 VDD.n1108 VDD.t1161 20.995
R7456 VDD.n1180 VDD.t1143 20.995
R7457 VDD.n1252 VDD.t1167 20.995
R7458 VDD.n1324 VDD.t1123 20.995
R7459 VDD.n1396 VDD.t1141 20.995
R7460 VDD.n1468 VDD.t1109 20.995
R7461 VDD.n1540 VDD.t1145 20.995
R7462 VDD.n1620 VDD.t1151 20.995
R7463 VDD.n537 VDD.t1147 20.995
R7464 VDD.n600 VDD.t1115 20.995
R7465 VDD.n597 VDD.t1125 20.628
R7466 VDD.n673 VDD.t1131 20.628
R7467 VDD.n745 VDD.t1105 20.628
R7468 VDD.n817 VDD.t1135 20.628
R7469 VDD.n889 VDD.t1107 20.628
R7470 VDD.n961 VDD.t1111 20.628
R7471 VDD.n1033 VDD.t1133 20.628
R7472 VDD.n1105 VDD.t1117 20.628
R7473 VDD.n1177 VDD.t1137 20.628
R7474 VDD.n1249 VDD.t1159 20.628
R7475 VDD.n1321 VDD.t1113 20.628
R7476 VDD.n1393 VDD.t1165 20.628
R7477 VDD.n1465 VDD.t1121 20.628
R7478 VDD.n1537 VDD.t1129 20.628
R7479 VDD.n1617 VDD.t1153 20.628
R7480 VDD.n534 VDD.t1155 20.628
R7481 VDD.n17 VDD.n16 19.954
R7482 VDD.n29 VDD.n28 19.954
R7483 VDD.n49 VDD.n48 19.954
R7484 VDD.n61 VDD.n60 19.954
R7485 VDD.n81 VDD.n80 19.954
R7486 VDD.n93 VDD.n92 19.954
R7487 VDD.n113 VDD.n112 19.954
R7488 VDD.n125 VDD.n124 19.954
R7489 VDD.n145 VDD.n144 19.954
R7490 VDD.n157 VDD.n156 19.954
R7491 VDD.n177 VDD.n176 19.954
R7492 VDD.n189 VDD.n188 19.954
R7493 VDD.n209 VDD.n208 19.954
R7494 VDD.n221 VDD.n220 19.954
R7495 VDD.n241 VDD.n240 19.954
R7496 VDD.n253 VDD.n252 19.954
R7497 VDD.n273 VDD.n272 19.954
R7498 VDD.n285 VDD.n284 19.954
R7499 VDD.n305 VDD.n304 19.954
R7500 VDD.n317 VDD.n316 19.954
R7501 VDD.n337 VDD.n336 19.954
R7502 VDD.n349 VDD.n348 19.954
R7503 VDD.n369 VDD.n368 19.954
R7504 VDD.n381 VDD.n380 19.954
R7505 VDD.n401 VDD.n400 19.954
R7506 VDD.n413 VDD.n412 19.954
R7507 VDD.n433 VDD.n432 19.954
R7508 VDD.n445 VDD.n444 19.954
R7509 VDD.n465 VDD.n464 19.954
R7510 VDD.n477 VDD.n476 19.954
R7511 VDD.n497 VDD.n496 19.954
R7512 VDD.n509 VDD.n508 19.954
R7513 VDD.n588 VDD.t2056 9.895
R7514 VDD.n660 VDD.t2022 9.895
R7515 VDD.n732 VDD.t2043 9.895
R7516 VDD.n804 VDD.t2083 9.895
R7517 VDD.n876 VDD.t2025 9.895
R7518 VDD.n948 VDD.t2088 9.895
R7519 VDD.n1020 VDD.t2087 9.895
R7520 VDD.n1092 VDD.t2075 9.895
R7521 VDD.n1164 VDD.t2017 9.895
R7522 VDD.n1236 VDD.t2055 9.895
R7523 VDD.n1308 VDD.t2080 9.895
R7524 VDD.n1380 VDD.t2042 9.895
R7525 VDD.n1452 VDD.t2084 9.895
R7526 VDD.n1524 VDD.t2048 9.895
R7527 VDD.n1596 VDD.t2074 9.895
R7528 VDD.n1607 VDD.t2065 9.895
R7529 VDD.n681 VDD.n680 8
R7530 VDD.n753 VDD.n752 8
R7531 VDD.n825 VDD.n824 8
R7532 VDD.n897 VDD.n896 8
R7533 VDD.n969 VDD.n968 8
R7534 VDD.n1041 VDD.n1040 8
R7535 VDD.n1113 VDD.n1112 8
R7536 VDD.n1185 VDD.n1184 8
R7537 VDD.n1257 VDD.n1256 8
R7538 VDD.n1329 VDD.n1328 8
R7539 VDD.n1401 VDD.n1400 8
R7540 VDD.n1473 VDD.n1472 8
R7541 VDD.n1545 VDD.n1544 8
R7542 VDD.n1625 VDD.n1624 8
R7543 VDD.n541 VDD.n540 8
R7544 VDD.n606 VDD.n605 8
R7545 VDD.n1678 VDD.n1677 7.566
R7546 VDD.n1623 VDD.n1622 6.744
R7547 VDD.n539 VDD.n538 6.436
R7548 VDD.n679 VDD.n678 6.405
R7549 VDD.n751 VDD.n750 6.405
R7550 VDD.n823 VDD.n822 6.405
R7551 VDD.n895 VDD.n894 6.405
R7552 VDD.n967 VDD.n966 6.405
R7553 VDD.n1039 VDD.n1038 6.405
R7554 VDD.n1111 VDD.n1110 6.405
R7555 VDD.n1183 VDD.n1182 6.405
R7556 VDD.n1255 VDD.n1254 6.405
R7557 VDD.n1327 VDD.n1326 6.405
R7558 VDD.n1399 VDD.n1398 6.405
R7559 VDD.n1471 VDD.n1470 6.405
R7560 VDD.n1543 VDD.n1542 6.405
R7561 VDD.n604 VDD.n603 6.405
R7562 VDD.n596 VDD.n595 6.065
R7563 VDD.n740 VDD.n739 6.065
R7564 VDD.n812 VDD.n811 6.065
R7565 VDD.n884 VDD.n883 6.065
R7566 VDD.n956 VDD.n955 6.065
R7567 VDD.n1028 VDD.n1027 6.065
R7568 VDD.n1100 VDD.n1099 6.065
R7569 VDD.n1172 VDD.n1171 6.065
R7570 VDD.n1244 VDD.n1243 6.065
R7571 VDD.n1316 VDD.n1315 6.065
R7572 VDD.n1388 VDD.n1387 6.065
R7573 VDD.n1460 VDD.n1459 6.065
R7574 VDD.n1532 VDD.n1531 6.065
R7575 VDD.n1604 VDD.n1603 6.065
R7576 VDD.n1676 VDD.n1606 6.065
R7577 VDD.n668 VDD.n667 6.065
R7578 VDD.n2 VDD.n1 4.574
R7579 VDD.n27 VDD.n26 4.574
R7580 VDD.n6 VDD.n5 4.574
R7581 VDD.n12 VDD.n11 4.574
R7582 VDD.n33 VDD.n32 4.574
R7583 VDD.n59 VDD.n58 4.574
R7584 VDD.n39 VDD.n38 4.574
R7585 VDD.n44 VDD.n43 4.574
R7586 VDD.n66 VDD.n65 4.574
R7587 VDD.n91 VDD.n90 4.574
R7588 VDD.n70 VDD.n69 4.574
R7589 VDD.n76 VDD.n75 4.574
R7590 VDD.n97 VDD.n96 4.574
R7591 VDD.n123 VDD.n122 4.574
R7592 VDD.n102 VDD.n101 4.574
R7593 VDD.n108 VDD.n107 4.574
R7594 VDD.n129 VDD.n128 4.574
R7595 VDD.n155 VDD.n154 4.574
R7596 VDD.n134 VDD.n133 4.574
R7597 VDD.n140 VDD.n139 4.574
R7598 VDD.n162 VDD.n161 4.574
R7599 VDD.n187 VDD.n186 4.574
R7600 VDD.n167 VDD.n166 4.574
R7601 VDD.n172 VDD.n171 4.574
R7602 VDD.n193 VDD.n192 4.574
R7603 VDD.n219 VDD.n218 4.574
R7604 VDD.n198 VDD.n197 4.574
R7605 VDD.n204 VDD.n203 4.574
R7606 VDD.n225 VDD.n224 4.574
R7607 VDD.n251 VDD.n250 4.574
R7608 VDD.n230 VDD.n229 4.574
R7609 VDD.n236 VDD.n235 4.574
R7610 VDD.n257 VDD.n256 4.574
R7611 VDD.n283 VDD.n282 4.574
R7612 VDD.n263 VDD.n262 4.574
R7613 VDD.n268 VDD.n267 4.574
R7614 VDD.n289 VDD.n288 4.574
R7615 VDD.n315 VDD.n314 4.574
R7616 VDD.n294 VDD.n293 4.574
R7617 VDD.n300 VDD.n299 4.574
R7618 VDD.n321 VDD.n320 4.574
R7619 VDD.n347 VDD.n346 4.574
R7620 VDD.n327 VDD.n326 4.574
R7621 VDD.n332 VDD.n331 4.574
R7622 VDD.n354 VDD.n353 4.574
R7623 VDD.n379 VDD.n378 4.574
R7624 VDD.n358 VDD.n357 4.574
R7625 VDD.n364 VDD.n363 4.574
R7626 VDD.n386 VDD.n385 4.574
R7627 VDD.n411 VDD.n410 4.574
R7628 VDD.n391 VDD.n390 4.574
R7629 VDD.n396 VDD.n395 4.574
R7630 VDD.n418 VDD.n417 4.574
R7631 VDD.n443 VDD.n442 4.574
R7632 VDD.n422 VDD.n421 4.574
R7633 VDD.n428 VDD.n427 4.574
R7634 VDD.n449 VDD.n448 4.574
R7635 VDD.n475 VDD.n474 4.574
R7636 VDD.n455 VDD.n454 4.574
R7637 VDD.n460 VDD.n459 4.574
R7638 VDD.n482 VDD.n481 4.574
R7639 VDD.n507 VDD.n506 4.574
R7640 VDD.n486 VDD.n485 4.574
R7641 VDD.n492 VDD.n491 4.574
R7642 VDD.n599 VDD.n598 4.574
R7643 VDD.n675 VDD.n674 4.574
R7644 VDD.n747 VDD.n746 4.574
R7645 VDD.n819 VDD.n818 4.574
R7646 VDD.n891 VDD.n890 4.574
R7647 VDD.n963 VDD.n962 4.574
R7648 VDD.n1035 VDD.n1034 4.574
R7649 VDD.n1107 VDD.n1106 4.574
R7650 VDD.n1179 VDD.n1178 4.574
R7651 VDD.n1251 VDD.n1250 4.574
R7652 VDD.n1323 VDD.n1322 4.574
R7653 VDD.n1395 VDD.n1394 4.574
R7654 VDD.n1467 VDD.n1466 4.574
R7655 VDD.n1539 VDD.n1538 4.574
R7656 VDD.n1619 VDD.n1618 4.574
R7657 VDD.n536 VDD.n535 4.574
R7658 VDD.n680 VDD.n679 4.5
R7659 VDD.n752 VDD.n751 4.5
R7660 VDD.n824 VDD.n823 4.5
R7661 VDD.n896 VDD.n895 4.5
R7662 VDD.n968 VDD.n967 4.5
R7663 VDD.n1040 VDD.n1039 4.5
R7664 VDD.n1112 VDD.n1111 4.5
R7665 VDD.n1184 VDD.n1183 4.5
R7666 VDD.n1256 VDD.n1255 4.5
R7667 VDD.n1328 VDD.n1327 4.5
R7668 VDD.n1400 VDD.n1399 4.5
R7669 VDD.n1472 VDD.n1471 4.5
R7670 VDD.n1544 VDD.n1543 4.5
R7671 VDD.n1624 VDD.n1623 4.5
R7672 VDD.n540 VDD.n539 4.5
R7673 VDD.n605 VDD.n604 4.5
R7674 VDD.n28 VDD.n27 4.491
R7675 VDD.n60 VDD.n59 4.491
R7676 VDD.n92 VDD.n91 4.491
R7677 VDD.n124 VDD.n123 4.491
R7678 VDD.n156 VDD.n155 4.491
R7679 VDD.n188 VDD.n187 4.491
R7680 VDD.n220 VDD.n219 4.491
R7681 VDD.n252 VDD.n251 4.491
R7682 VDD.n284 VDD.n283 4.491
R7683 VDD.n316 VDD.n315 4.491
R7684 VDD.n348 VDD.n347 4.491
R7685 VDD.n380 VDD.n379 4.491
R7686 VDD.n412 VDD.n411 4.491
R7687 VDD.n444 VDD.n443 4.491
R7688 VDD.n476 VDD.n475 4.491
R7689 VDD.n508 VDD.n507 4.491
R7690 VDD.n18 VDD.n9 4.49
R7691 VDD.n18 VDD.n7 4.49
R7692 VDD.n30 VDD.n4 4.49
R7693 VDD.n30 VDD.n0 4.49
R7694 VDD.n50 VDD.n41 4.49
R7695 VDD.n50 VDD.n37 4.49
R7696 VDD.n62 VDD.n36 4.49
R7697 VDD.n62 VDD.n34 4.49
R7698 VDD.n82 VDD.n73 4.49
R7699 VDD.n82 VDD.n71 4.49
R7700 VDD.n94 VDD.n68 4.49
R7701 VDD.n94 VDD.n64 4.49
R7702 VDD.n114 VDD.n105 4.49
R7703 VDD.n114 VDD.n103 4.49
R7704 VDD.n126 VDD.n100 4.49
R7705 VDD.n126 VDD.n98 4.49
R7706 VDD.n146 VDD.n137 4.49
R7707 VDD.n146 VDD.n135 4.49
R7708 VDD.n158 VDD.n132 4.49
R7709 VDD.n158 VDD.n130 4.49
R7710 VDD.n178 VDD.n169 4.49
R7711 VDD.n178 VDD.n165 4.49
R7712 VDD.n190 VDD.n164 4.49
R7713 VDD.n190 VDD.n160 4.49
R7714 VDD.n210 VDD.n201 4.49
R7715 VDD.n210 VDD.n199 4.49
R7716 VDD.n222 VDD.n196 4.49
R7717 VDD.n222 VDD.n194 4.49
R7718 VDD.n242 VDD.n233 4.49
R7719 VDD.n242 VDD.n231 4.49
R7720 VDD.n254 VDD.n228 4.49
R7721 VDD.n254 VDD.n226 4.49
R7722 VDD.n274 VDD.n265 4.49
R7723 VDD.n274 VDD.n261 4.49
R7724 VDD.n286 VDD.n260 4.49
R7725 VDD.n286 VDD.n258 4.49
R7726 VDD.n306 VDD.n297 4.49
R7727 VDD.n306 VDD.n295 4.49
R7728 VDD.n318 VDD.n292 4.49
R7729 VDD.n318 VDD.n290 4.49
R7730 VDD.n338 VDD.n329 4.49
R7731 VDD.n338 VDD.n325 4.49
R7732 VDD.n350 VDD.n324 4.49
R7733 VDD.n350 VDD.n322 4.49
R7734 VDD.n370 VDD.n361 4.49
R7735 VDD.n370 VDD.n359 4.49
R7736 VDD.n382 VDD.n356 4.49
R7737 VDD.n382 VDD.n352 4.49
R7738 VDD.n402 VDD.n393 4.49
R7739 VDD.n402 VDD.n389 4.49
R7740 VDD.n414 VDD.n388 4.49
R7741 VDD.n414 VDD.n384 4.49
R7742 VDD.n434 VDD.n425 4.49
R7743 VDD.n434 VDD.n423 4.49
R7744 VDD.n446 VDD.n420 4.49
R7745 VDD.n446 VDD.n416 4.49
R7746 VDD.n466 VDD.n457 4.49
R7747 VDD.n466 VDD.n453 4.49
R7748 VDD.n478 VDD.n452 4.49
R7749 VDD.n478 VDD.n450 4.49
R7750 VDD.n498 VDD.n489 4.49
R7751 VDD.n498 VDD.n487 4.49
R7752 VDD.n510 VDD.n484 4.49
R7753 VDD.n510 VDD.n480 4.49
R7754 VDD.n735 VDD.n734 4.207
R7755 VDD.n807 VDD.n806 4.207
R7756 VDD.n879 VDD.n878 4.207
R7757 VDD.n951 VDD.n950 4.207
R7758 VDD.n1023 VDD.n1022 4.207
R7759 VDD.n1095 VDD.n1094 4.207
R7760 VDD.n1167 VDD.n1166 4.207
R7761 VDD.n1239 VDD.n1238 4.207
R7762 VDD.n1311 VDD.n1310 4.207
R7763 VDD.n1383 VDD.n1382 4.207
R7764 VDD.n1455 VDD.n1454 4.207
R7765 VDD.n1527 VDD.n1526 4.207
R7766 VDD.n1599 VDD.n1598 4.207
R7767 VDD.n663 VDD.n662 4.207
R7768 VDD.n702 VDD.n701 4.206
R7769 VDD.n720 VDD.n719 4.206
R7770 VDD.n688 VDD.n672 4.206
R7771 VDD.n774 VDD.n773 4.206
R7772 VDD.n792 VDD.n791 4.206
R7773 VDD.n760 VDD.n744 4.206
R7774 VDD.n846 VDD.n845 4.206
R7775 VDD.n864 VDD.n863 4.206
R7776 VDD.n832 VDD.n816 4.206
R7777 VDD.n918 VDD.n917 4.206
R7778 VDD.n936 VDD.n935 4.206
R7779 VDD.n904 VDD.n888 4.206
R7780 VDD.n990 VDD.n989 4.206
R7781 VDD.n1008 VDD.n1007 4.206
R7782 VDD.n976 VDD.n960 4.206
R7783 VDD.n1062 VDD.n1061 4.206
R7784 VDD.n1080 VDD.n1079 4.206
R7785 VDD.n1048 VDD.n1032 4.206
R7786 VDD.n1134 VDD.n1133 4.206
R7787 VDD.n1152 VDD.n1151 4.206
R7788 VDD.n1120 VDD.n1104 4.206
R7789 VDD.n1206 VDD.n1205 4.206
R7790 VDD.n1224 VDD.n1223 4.206
R7791 VDD.n1192 VDD.n1176 4.206
R7792 VDD.n1278 VDD.n1277 4.206
R7793 VDD.n1296 VDD.n1295 4.206
R7794 VDD.n1264 VDD.n1248 4.206
R7795 VDD.n1350 VDD.n1349 4.206
R7796 VDD.n1368 VDD.n1367 4.206
R7797 VDD.n1336 VDD.n1320 4.206
R7798 VDD.n1422 VDD.n1421 4.206
R7799 VDD.n1440 VDD.n1439 4.206
R7800 VDD.n1408 VDD.n1392 4.206
R7801 VDD.n1494 VDD.n1493 4.206
R7802 VDD.n1512 VDD.n1511 4.206
R7803 VDD.n1480 VDD.n1464 4.206
R7804 VDD.n1566 VDD.n1565 4.206
R7805 VDD.n1584 VDD.n1583 4.206
R7806 VDD.n1552 VDD.n1536 4.206
R7807 VDD.n1672 VDD.n1609 4.206
R7808 VDD.n1660 VDD.n1611 4.206
R7809 VDD.n1644 VDD.n1613 4.206
R7810 VDD.n1632 VDD.n1616 4.206
R7811 VDD.n576 VDD.n528 4.206
R7812 VDD.n560 VDD.n530 4.206
R7813 VDD.n548 VDD.n533 4.206
R7814 VDD.n616 VDD.n615 4.206
R7815 VDD.n630 VDD.n629 4.206
R7816 VDD.n648 VDD.n647 4.206
R7817 VDD.n591 VDD.n590 4.206
R7818 VDD.n20 VDD.n19 3.975
R7819 VDD.n52 VDD.n51 3.975
R7820 VDD.n84 VDD.n83 3.975
R7821 VDD.n116 VDD.n115 3.975
R7822 VDD.n148 VDD.n147 3.975
R7823 VDD.n180 VDD.n179 3.975
R7824 VDD.n212 VDD.n211 3.975
R7825 VDD.n244 VDD.n243 3.975
R7826 VDD.n276 VDD.n275 3.975
R7827 VDD.n308 VDD.n307 3.975
R7828 VDD.n340 VDD.n339 3.975
R7829 VDD.n372 VDD.n371 3.975
R7830 VDD.n404 VDD.n403 3.975
R7831 VDD.n436 VDD.n435 3.975
R7832 VDD.n468 VDD.n467 3.975
R7833 VDD.n500 VDD.n499 3.975
R7834 VDD.n512 VDD.n511 3.761
R7835 VDD.n15 VDD.n14 2.996
R7836 VDD.n47 VDD.n46 2.996
R7837 VDD.n79 VDD.n78 2.996
R7838 VDD.n111 VDD.n110 2.996
R7839 VDD.n143 VDD.n142 2.996
R7840 VDD.n175 VDD.n174 2.996
R7841 VDD.n207 VDD.n206 2.996
R7842 VDD.n239 VDD.n238 2.996
R7843 VDD.n271 VDD.n270 2.996
R7844 VDD.n303 VDD.n302 2.996
R7845 VDD.n335 VDD.n334 2.996
R7846 VDD.n367 VDD.n366 2.996
R7847 VDD.n399 VDD.n398 2.996
R7848 VDD.n431 VDD.n430 2.996
R7849 VDD.n463 VDD.n462 2.996
R7850 VDD.n495 VDD.n494 2.996
R7851 VDD.n682 VDD.n676 2.991
R7852 VDD.n754 VDD.n748 2.991
R7853 VDD.n826 VDD.n820 2.991
R7854 VDD.n898 VDD.n892 2.991
R7855 VDD.n970 VDD.n964 2.991
R7856 VDD.n1042 VDD.n1036 2.991
R7857 VDD.n1114 VDD.n1108 2.991
R7858 VDD.n1186 VDD.n1180 2.991
R7859 VDD.n1258 VDD.n1252 2.991
R7860 VDD.n1330 VDD.n1324 2.991
R7861 VDD.n1402 VDD.n1396 2.991
R7862 VDD.n1474 VDD.n1468 2.991
R7863 VDD.n1546 VDD.n1540 2.991
R7864 VDD.n1626 VDD.n1620 2.991
R7865 VDD.n542 VDD.n537 2.991
R7866 VDD.n607 VDD.n600 2.991
R7867 VDD.n524 VDD.n95 2.396
R7868 VDD.n513 VDD.n447 2.396
R7869 VDD.n526 VDD.n31 2.387
R7870 VDD.n525 VDD.n63 2.387
R7871 VDD.n519 VDD.n255 2.387
R7872 VDD.n516 VDD.n351 2.378
R7873 VDD.n512 VDD.n479 2.378
R7874 VDD.n522 VDD.n159 2.369
R7875 VDD.n515 VDD.n383 2.369
R7876 VDD.n521 VDD.n191 2.36
R7877 VDD.n520 VDD.n223 2.36
R7878 VDD.n518 VDD.n287 2.36
R7879 VDD.n517 VDD.n319 2.36
R7880 VDD.n514 VDD.n415 2.36
R7881 VDD.n523 VDD.n127 2.352
R7882 VDD.n513 VDD.n512 1.849
R7883 VDD.n514 VDD.n513 1.849
R7884 VDD.n515 VDD.n514 1.844
R7885 VDD.n516 VDD.n515 1.844
R7886 VDD.n517 VDD.n516 1.841
R7887 VDD.n518 VDD.n517 1.841
R7888 VDD.n519 VDD.n518 1.841
R7889 VDD.n520 VDD.n519 1.841
R7890 VDD.n521 VDD.n520 1.841
R7891 VDD.n522 VDD.n521 1.841
R7892 VDD.n525 VDD.n524 1.841
R7893 VDD.n523 VDD.n522 1.838
R7894 VDD.n524 VDD.n523 1.838
R7895 VDD.n526 VDD.n525 1.791
R7896 VDD.n669 VDD.n596 1.561
R7897 VDD.n14 VDD.n13 1.41
R7898 VDD.n46 VDD.n45 1.41
R7899 VDD.n78 VDD.n77 1.41
R7900 VDD.n110 VDD.n109 1.41
R7901 VDD.n142 VDD.n141 1.41
R7902 VDD.n174 VDD.n173 1.41
R7903 VDD.n206 VDD.n205 1.41
R7904 VDD.n238 VDD.n237 1.41
R7905 VDD.n270 VDD.n269 1.41
R7906 VDD.n302 VDD.n301 1.41
R7907 VDD.n334 VDD.n333 1.41
R7908 VDD.n366 VDD.n365 1.41
R7909 VDD.n398 VDD.n397 1.41
R7910 VDD.n430 VDD.n429 1.41
R7911 VDD.n462 VDD.n461 1.41
R7912 VDD.n494 VDD.n493 1.41
R7913 VDD.n4 VDD.n3 1.402
R7914 VDD.n24 VDD.n23 1.402
R7915 VDD.n9 VDD.n8 1.402
R7916 VDD.n36 VDD.n35 1.402
R7917 VDD.n56 VDD.n55 1.402
R7918 VDD.n41 VDD.n40 1.402
R7919 VDD.n68 VDD.n67 1.402
R7920 VDD.n88 VDD.n87 1.402
R7921 VDD.n73 VDD.n72 1.402
R7922 VDD.n100 VDD.n99 1.402
R7923 VDD.n120 VDD.n119 1.402
R7924 VDD.n105 VDD.n104 1.402
R7925 VDD.n132 VDD.n131 1.402
R7926 VDD.n152 VDD.n151 1.402
R7927 VDD.n137 VDD.n136 1.402
R7928 VDD.n164 VDD.n163 1.402
R7929 VDD.n184 VDD.n183 1.402
R7930 VDD.n169 VDD.n168 1.402
R7931 VDD.n196 VDD.n195 1.402
R7932 VDD.n216 VDD.n215 1.402
R7933 VDD.n201 VDD.n200 1.402
R7934 VDD.n228 VDD.n227 1.402
R7935 VDD.n248 VDD.n247 1.402
R7936 VDD.n233 VDD.n232 1.402
R7937 VDD.n260 VDD.n259 1.402
R7938 VDD.n280 VDD.n279 1.402
R7939 VDD.n265 VDD.n264 1.402
R7940 VDD.n292 VDD.n291 1.402
R7941 VDD.n312 VDD.n311 1.402
R7942 VDD.n297 VDD.n296 1.402
R7943 VDD.n324 VDD.n323 1.402
R7944 VDD.n344 VDD.n343 1.402
R7945 VDD.n329 VDD.n328 1.402
R7946 VDD.n356 VDD.n355 1.402
R7947 VDD.n376 VDD.n375 1.402
R7948 VDD.n361 VDD.n360 1.402
R7949 VDD.n388 VDD.n387 1.402
R7950 VDD.n408 VDD.n407 1.402
R7951 VDD.n393 VDD.n392 1.402
R7952 VDD.n420 VDD.n419 1.402
R7953 VDD.n440 VDD.n439 1.402
R7954 VDD.n425 VDD.n424 1.402
R7955 VDD.n452 VDD.n451 1.402
R7956 VDD.n472 VDD.n471 1.402
R7957 VDD.n457 VDD.n456 1.402
R7958 VDD.n484 VDD.n483 1.402
R7959 VDD.n504 VDD.n503 1.402
R7960 VDD.n489 VDD.n488 1.402
R7961 VDD.n684 VDD.n683 1.367
R7962 VDD.n756 VDD.n755 1.367
R7963 VDD.n828 VDD.n827 1.367
R7964 VDD.n900 VDD.n899 1.367
R7965 VDD.n972 VDD.n971 1.367
R7966 VDD.n1044 VDD.n1043 1.367
R7967 VDD.n1116 VDD.n1115 1.367
R7968 VDD.n1188 VDD.n1187 1.367
R7969 VDD.n1260 VDD.n1259 1.367
R7970 VDD.n1332 VDD.n1331 1.367
R7971 VDD.n1404 VDD.n1403 1.367
R7972 VDD.n1476 VDD.n1475 1.367
R7973 VDD.n1548 VDD.n1547 1.367
R7974 VDD.n1628 VDD.n1627 1.367
R7975 VDD.n544 VDD.n543 1.367
R7976 VDD.n609 VDD.n608 1.367
R7977 VDD.n689 VDD.n688 1.133
R7978 VDD.n691 VDD.n690 1.133
R7979 VDD.n693 VDD.n692 1.133
R7980 VDD.n695 VDD.n694 1.133
R7981 VDD.n697 VDD.n696 1.133
R7982 VDD.n699 VDD.n698 1.133
R7983 VDD.n703 VDD.n702 1.133
R7984 VDD.n705 VDD.n704 1.133
R7985 VDD.n707 VDD.n706 1.133
R7986 VDD.n709 VDD.n708 1.133
R7987 VDD.n711 VDD.n710 1.133
R7988 VDD.n713 VDD.n712 1.133
R7989 VDD.n715 VDD.n714 1.133
R7990 VDD.n717 VDD.n716 1.133
R7991 VDD.n721 VDD.n720 1.133
R7992 VDD.n723 VDD.n722 1.133
R7993 VDD.n725 VDD.n724 1.133
R7994 VDD.n727 VDD.n726 1.133
R7995 VDD.n729 VDD.n728 1.133
R7996 VDD.n731 VDD.n730 1.133
R7997 VDD.n738 VDD.n737 1.133
R7998 VDD.n736 VDD.n735 1.133
R7999 VDD.n687 VDD.n686 1.133
R8000 VDD.n685 VDD.n684 1.133
R8001 VDD.n761 VDD.n760 1.133
R8002 VDD.n763 VDD.n762 1.133
R8003 VDD.n765 VDD.n764 1.133
R8004 VDD.n767 VDD.n766 1.133
R8005 VDD.n769 VDD.n768 1.133
R8006 VDD.n771 VDD.n770 1.133
R8007 VDD.n775 VDD.n774 1.133
R8008 VDD.n777 VDD.n776 1.133
R8009 VDD.n779 VDD.n778 1.133
R8010 VDD.n781 VDD.n780 1.133
R8011 VDD.n783 VDD.n782 1.133
R8012 VDD.n785 VDD.n784 1.133
R8013 VDD.n787 VDD.n786 1.133
R8014 VDD.n789 VDD.n788 1.133
R8015 VDD.n793 VDD.n792 1.133
R8016 VDD.n795 VDD.n794 1.133
R8017 VDD.n797 VDD.n796 1.133
R8018 VDD.n799 VDD.n798 1.133
R8019 VDD.n801 VDD.n800 1.133
R8020 VDD.n803 VDD.n802 1.133
R8021 VDD.n810 VDD.n809 1.133
R8022 VDD.n808 VDD.n807 1.133
R8023 VDD.n759 VDD.n758 1.133
R8024 VDD.n757 VDD.n756 1.133
R8025 VDD.n833 VDD.n832 1.133
R8026 VDD.n835 VDD.n834 1.133
R8027 VDD.n837 VDD.n836 1.133
R8028 VDD.n839 VDD.n838 1.133
R8029 VDD.n841 VDD.n840 1.133
R8030 VDD.n843 VDD.n842 1.133
R8031 VDD.n847 VDD.n846 1.133
R8032 VDD.n849 VDD.n848 1.133
R8033 VDD.n851 VDD.n850 1.133
R8034 VDD.n853 VDD.n852 1.133
R8035 VDD.n855 VDD.n854 1.133
R8036 VDD.n857 VDD.n856 1.133
R8037 VDD.n859 VDD.n858 1.133
R8038 VDD.n861 VDD.n860 1.133
R8039 VDD.n865 VDD.n864 1.133
R8040 VDD.n867 VDD.n866 1.133
R8041 VDD.n869 VDD.n868 1.133
R8042 VDD.n871 VDD.n870 1.133
R8043 VDD.n873 VDD.n872 1.133
R8044 VDD.n875 VDD.n874 1.133
R8045 VDD.n882 VDD.n881 1.133
R8046 VDD.n880 VDD.n879 1.133
R8047 VDD.n831 VDD.n830 1.133
R8048 VDD.n829 VDD.n828 1.133
R8049 VDD.n905 VDD.n904 1.133
R8050 VDD.n907 VDD.n906 1.133
R8051 VDD.n909 VDD.n908 1.133
R8052 VDD.n911 VDD.n910 1.133
R8053 VDD.n913 VDD.n912 1.133
R8054 VDD.n915 VDD.n914 1.133
R8055 VDD.n919 VDD.n918 1.133
R8056 VDD.n921 VDD.n920 1.133
R8057 VDD.n923 VDD.n922 1.133
R8058 VDD.n925 VDD.n924 1.133
R8059 VDD.n927 VDD.n926 1.133
R8060 VDD.n929 VDD.n928 1.133
R8061 VDD.n931 VDD.n930 1.133
R8062 VDD.n933 VDD.n932 1.133
R8063 VDD.n937 VDD.n936 1.133
R8064 VDD.n939 VDD.n938 1.133
R8065 VDD.n941 VDD.n940 1.133
R8066 VDD.n943 VDD.n942 1.133
R8067 VDD.n945 VDD.n944 1.133
R8068 VDD.n947 VDD.n946 1.133
R8069 VDD.n954 VDD.n953 1.133
R8070 VDD.n952 VDD.n951 1.133
R8071 VDD.n903 VDD.n902 1.133
R8072 VDD.n901 VDD.n900 1.133
R8073 VDD.n977 VDD.n976 1.133
R8074 VDD.n979 VDD.n978 1.133
R8075 VDD.n981 VDD.n980 1.133
R8076 VDD.n983 VDD.n982 1.133
R8077 VDD.n985 VDD.n984 1.133
R8078 VDD.n987 VDD.n986 1.133
R8079 VDD.n991 VDD.n990 1.133
R8080 VDD.n993 VDD.n992 1.133
R8081 VDD.n995 VDD.n994 1.133
R8082 VDD.n997 VDD.n996 1.133
R8083 VDD.n999 VDD.n998 1.133
R8084 VDD.n1001 VDD.n1000 1.133
R8085 VDD.n1003 VDD.n1002 1.133
R8086 VDD.n1005 VDD.n1004 1.133
R8087 VDD.n1009 VDD.n1008 1.133
R8088 VDD.n1011 VDD.n1010 1.133
R8089 VDD.n1013 VDD.n1012 1.133
R8090 VDD.n1015 VDD.n1014 1.133
R8091 VDD.n1017 VDD.n1016 1.133
R8092 VDD.n1019 VDD.n1018 1.133
R8093 VDD.n1026 VDD.n1025 1.133
R8094 VDD.n1024 VDD.n1023 1.133
R8095 VDD.n975 VDD.n974 1.133
R8096 VDD.n973 VDD.n972 1.133
R8097 VDD.n1049 VDD.n1048 1.133
R8098 VDD.n1051 VDD.n1050 1.133
R8099 VDD.n1053 VDD.n1052 1.133
R8100 VDD.n1055 VDD.n1054 1.133
R8101 VDD.n1057 VDD.n1056 1.133
R8102 VDD.n1059 VDD.n1058 1.133
R8103 VDD.n1063 VDD.n1062 1.133
R8104 VDD.n1065 VDD.n1064 1.133
R8105 VDD.n1067 VDD.n1066 1.133
R8106 VDD.n1069 VDD.n1068 1.133
R8107 VDD.n1071 VDD.n1070 1.133
R8108 VDD.n1073 VDD.n1072 1.133
R8109 VDD.n1075 VDD.n1074 1.133
R8110 VDD.n1077 VDD.n1076 1.133
R8111 VDD.n1081 VDD.n1080 1.133
R8112 VDD.n1083 VDD.n1082 1.133
R8113 VDD.n1085 VDD.n1084 1.133
R8114 VDD.n1087 VDD.n1086 1.133
R8115 VDD.n1089 VDD.n1088 1.133
R8116 VDD.n1091 VDD.n1090 1.133
R8117 VDD.n1098 VDD.n1097 1.133
R8118 VDD.n1096 VDD.n1095 1.133
R8119 VDD.n1047 VDD.n1046 1.133
R8120 VDD.n1045 VDD.n1044 1.133
R8121 VDD.n1121 VDD.n1120 1.133
R8122 VDD.n1123 VDD.n1122 1.133
R8123 VDD.n1125 VDD.n1124 1.133
R8124 VDD.n1127 VDD.n1126 1.133
R8125 VDD.n1129 VDD.n1128 1.133
R8126 VDD.n1131 VDD.n1130 1.133
R8127 VDD.n1135 VDD.n1134 1.133
R8128 VDD.n1137 VDD.n1136 1.133
R8129 VDD.n1139 VDD.n1138 1.133
R8130 VDD.n1141 VDD.n1140 1.133
R8131 VDD.n1143 VDD.n1142 1.133
R8132 VDD.n1145 VDD.n1144 1.133
R8133 VDD.n1147 VDD.n1146 1.133
R8134 VDD.n1149 VDD.n1148 1.133
R8135 VDD.n1153 VDD.n1152 1.133
R8136 VDD.n1155 VDD.n1154 1.133
R8137 VDD.n1157 VDD.n1156 1.133
R8138 VDD.n1159 VDD.n1158 1.133
R8139 VDD.n1161 VDD.n1160 1.133
R8140 VDD.n1163 VDD.n1162 1.133
R8141 VDD.n1170 VDD.n1169 1.133
R8142 VDD.n1168 VDD.n1167 1.133
R8143 VDD.n1119 VDD.n1118 1.133
R8144 VDD.n1117 VDD.n1116 1.133
R8145 VDD.n1193 VDD.n1192 1.133
R8146 VDD.n1195 VDD.n1194 1.133
R8147 VDD.n1197 VDD.n1196 1.133
R8148 VDD.n1199 VDD.n1198 1.133
R8149 VDD.n1201 VDD.n1200 1.133
R8150 VDD.n1203 VDD.n1202 1.133
R8151 VDD.n1207 VDD.n1206 1.133
R8152 VDD.n1209 VDD.n1208 1.133
R8153 VDD.n1211 VDD.n1210 1.133
R8154 VDD.n1213 VDD.n1212 1.133
R8155 VDD.n1215 VDD.n1214 1.133
R8156 VDD.n1217 VDD.n1216 1.133
R8157 VDD.n1219 VDD.n1218 1.133
R8158 VDD.n1221 VDD.n1220 1.133
R8159 VDD.n1225 VDD.n1224 1.133
R8160 VDD.n1227 VDD.n1226 1.133
R8161 VDD.n1229 VDD.n1228 1.133
R8162 VDD.n1231 VDD.n1230 1.133
R8163 VDD.n1233 VDD.n1232 1.133
R8164 VDD.n1235 VDD.n1234 1.133
R8165 VDD.n1242 VDD.n1241 1.133
R8166 VDD.n1240 VDD.n1239 1.133
R8167 VDD.n1191 VDD.n1190 1.133
R8168 VDD.n1189 VDD.n1188 1.133
R8169 VDD.n1265 VDD.n1264 1.133
R8170 VDD.n1267 VDD.n1266 1.133
R8171 VDD.n1269 VDD.n1268 1.133
R8172 VDD.n1271 VDD.n1270 1.133
R8173 VDD.n1273 VDD.n1272 1.133
R8174 VDD.n1275 VDD.n1274 1.133
R8175 VDD.n1279 VDD.n1278 1.133
R8176 VDD.n1281 VDD.n1280 1.133
R8177 VDD.n1283 VDD.n1282 1.133
R8178 VDD.n1285 VDD.n1284 1.133
R8179 VDD.n1287 VDD.n1286 1.133
R8180 VDD.n1289 VDD.n1288 1.133
R8181 VDD.n1291 VDD.n1290 1.133
R8182 VDD.n1293 VDD.n1292 1.133
R8183 VDD.n1297 VDD.n1296 1.133
R8184 VDD.n1299 VDD.n1298 1.133
R8185 VDD.n1301 VDD.n1300 1.133
R8186 VDD.n1303 VDD.n1302 1.133
R8187 VDD.n1305 VDD.n1304 1.133
R8188 VDD.n1307 VDD.n1306 1.133
R8189 VDD.n1314 VDD.n1313 1.133
R8190 VDD.n1312 VDD.n1311 1.133
R8191 VDD.n1263 VDD.n1262 1.133
R8192 VDD.n1261 VDD.n1260 1.133
R8193 VDD.n1337 VDD.n1336 1.133
R8194 VDD.n1339 VDD.n1338 1.133
R8195 VDD.n1341 VDD.n1340 1.133
R8196 VDD.n1343 VDD.n1342 1.133
R8197 VDD.n1345 VDD.n1344 1.133
R8198 VDD.n1347 VDD.n1346 1.133
R8199 VDD.n1351 VDD.n1350 1.133
R8200 VDD.n1353 VDD.n1352 1.133
R8201 VDD.n1355 VDD.n1354 1.133
R8202 VDD.n1357 VDD.n1356 1.133
R8203 VDD.n1359 VDD.n1358 1.133
R8204 VDD.n1361 VDD.n1360 1.133
R8205 VDD.n1363 VDD.n1362 1.133
R8206 VDD.n1365 VDD.n1364 1.133
R8207 VDD.n1369 VDD.n1368 1.133
R8208 VDD.n1371 VDD.n1370 1.133
R8209 VDD.n1373 VDD.n1372 1.133
R8210 VDD.n1375 VDD.n1374 1.133
R8211 VDD.n1377 VDD.n1376 1.133
R8212 VDD.n1379 VDD.n1378 1.133
R8213 VDD.n1386 VDD.n1385 1.133
R8214 VDD.n1384 VDD.n1383 1.133
R8215 VDD.n1335 VDD.n1334 1.133
R8216 VDD.n1333 VDD.n1332 1.133
R8217 VDD.n1409 VDD.n1408 1.133
R8218 VDD.n1411 VDD.n1410 1.133
R8219 VDD.n1413 VDD.n1412 1.133
R8220 VDD.n1415 VDD.n1414 1.133
R8221 VDD.n1417 VDD.n1416 1.133
R8222 VDD.n1419 VDD.n1418 1.133
R8223 VDD.n1423 VDD.n1422 1.133
R8224 VDD.n1425 VDD.n1424 1.133
R8225 VDD.n1427 VDD.n1426 1.133
R8226 VDD.n1429 VDD.n1428 1.133
R8227 VDD.n1431 VDD.n1430 1.133
R8228 VDD.n1433 VDD.n1432 1.133
R8229 VDD.n1435 VDD.n1434 1.133
R8230 VDD.n1437 VDD.n1436 1.133
R8231 VDD.n1441 VDD.n1440 1.133
R8232 VDD.n1443 VDD.n1442 1.133
R8233 VDD.n1445 VDD.n1444 1.133
R8234 VDD.n1447 VDD.n1446 1.133
R8235 VDD.n1449 VDD.n1448 1.133
R8236 VDD.n1451 VDD.n1450 1.133
R8237 VDD.n1458 VDD.n1457 1.133
R8238 VDD.n1456 VDD.n1455 1.133
R8239 VDD.n1407 VDD.n1406 1.133
R8240 VDD.n1405 VDD.n1404 1.133
R8241 VDD.n1481 VDD.n1480 1.133
R8242 VDD.n1483 VDD.n1482 1.133
R8243 VDD.n1485 VDD.n1484 1.133
R8244 VDD.n1487 VDD.n1486 1.133
R8245 VDD.n1489 VDD.n1488 1.133
R8246 VDD.n1491 VDD.n1490 1.133
R8247 VDD.n1495 VDD.n1494 1.133
R8248 VDD.n1497 VDD.n1496 1.133
R8249 VDD.n1499 VDD.n1498 1.133
R8250 VDD.n1501 VDD.n1500 1.133
R8251 VDD.n1503 VDD.n1502 1.133
R8252 VDD.n1505 VDD.n1504 1.133
R8253 VDD.n1507 VDD.n1506 1.133
R8254 VDD.n1509 VDD.n1508 1.133
R8255 VDD.n1513 VDD.n1512 1.133
R8256 VDD.n1515 VDD.n1514 1.133
R8257 VDD.n1517 VDD.n1516 1.133
R8258 VDD.n1519 VDD.n1518 1.133
R8259 VDD.n1521 VDD.n1520 1.133
R8260 VDD.n1523 VDD.n1522 1.133
R8261 VDD.n1530 VDD.n1529 1.133
R8262 VDD.n1528 VDD.n1527 1.133
R8263 VDD.n1479 VDD.n1478 1.133
R8264 VDD.n1477 VDD.n1476 1.133
R8265 VDD.n1553 VDD.n1552 1.133
R8266 VDD.n1555 VDD.n1554 1.133
R8267 VDD.n1557 VDD.n1556 1.133
R8268 VDD.n1559 VDD.n1558 1.133
R8269 VDD.n1561 VDD.n1560 1.133
R8270 VDD.n1563 VDD.n1562 1.133
R8271 VDD.n1567 VDD.n1566 1.133
R8272 VDD.n1569 VDD.n1568 1.133
R8273 VDD.n1571 VDD.n1570 1.133
R8274 VDD.n1573 VDD.n1572 1.133
R8275 VDD.n1575 VDD.n1574 1.133
R8276 VDD.n1577 VDD.n1576 1.133
R8277 VDD.n1579 VDD.n1578 1.133
R8278 VDD.n1581 VDD.n1580 1.133
R8279 VDD.n1585 VDD.n1584 1.133
R8280 VDD.n1587 VDD.n1586 1.133
R8281 VDD.n1589 VDD.n1588 1.133
R8282 VDD.n1591 VDD.n1590 1.133
R8283 VDD.n1593 VDD.n1592 1.133
R8284 VDD.n1595 VDD.n1594 1.133
R8285 VDD.n1602 VDD.n1601 1.133
R8286 VDD.n1600 VDD.n1599 1.133
R8287 VDD.n1551 VDD.n1550 1.133
R8288 VDD.n1549 VDD.n1548 1.133
R8289 VDD.n1675 VDD.n1674 1.133
R8290 VDD.n1673 VDD.n1672 1.133
R8291 VDD.n1671 VDD.n1670 1.133
R8292 VDD.n1669 VDD.n1668 1.133
R8293 VDD.n1667 VDD.n1666 1.133
R8294 VDD.n1665 VDD.n1664 1.133
R8295 VDD.n1663 VDD.n1662 1.133
R8296 VDD.n1661 VDD.n1660 1.133
R8297 VDD.n1659 VDD.n1658 1.133
R8298 VDD.n1657 VDD.n1656 1.133
R8299 VDD.n1655 VDD.n1654 1.133
R8300 VDD.n1653 VDD.n1652 1.133
R8301 VDD.n1651 VDD.n1650 1.133
R8302 VDD.n1649 VDD.n1648 1.133
R8303 VDD.n1647 VDD.n1646 1.133
R8304 VDD.n1645 VDD.n1644 1.133
R8305 VDD.n1643 VDD.n1642 1.133
R8306 VDD.n1641 VDD.n1640 1.133
R8307 VDD.n1639 VDD.n1638 1.133
R8308 VDD.n1637 VDD.n1636 1.133
R8309 VDD.n1635 VDD.n1634 1.133
R8310 VDD.n1633 VDD.n1632 1.133
R8311 VDD.n1631 VDD.n1630 1.133
R8312 VDD.n1629 VDD.n1628 1.133
R8313 VDD.n587 VDD.n586 1.133
R8314 VDD.n585 VDD.n584 1.133
R8315 VDD.n583 VDD.n582 1.133
R8316 VDD.n581 VDD.n580 1.133
R8317 VDD.n579 VDD.n578 1.133
R8318 VDD.n577 VDD.n576 1.133
R8319 VDD.n575 VDD.n574 1.133
R8320 VDD.n573 VDD.n572 1.133
R8321 VDD.n571 VDD.n570 1.133
R8322 VDD.n569 VDD.n568 1.133
R8323 VDD.n567 VDD.n566 1.133
R8324 VDD.n565 VDD.n564 1.133
R8325 VDD.n563 VDD.n562 1.133
R8326 VDD.n561 VDD.n560 1.133
R8327 VDD.n559 VDD.n558 1.133
R8328 VDD.n557 VDD.n556 1.133
R8329 VDD.n555 VDD.n554 1.133
R8330 VDD.n553 VDD.n552 1.133
R8331 VDD.n551 VDD.n550 1.133
R8332 VDD.n549 VDD.n548 1.133
R8333 VDD.n547 VDD.n546 1.133
R8334 VDD.n545 VDD.n544 1.133
R8335 VDD.n610 VDD.n609 1.133
R8336 VDD.n612 VDD.n611 1.133
R8337 VDD.n617 VDD.n616 1.133
R8338 VDD.n619 VDD.n618 1.133
R8339 VDD.n621 VDD.n620 1.133
R8340 VDD.n623 VDD.n622 1.133
R8341 VDD.n625 VDD.n624 1.133
R8342 VDD.n627 VDD.n626 1.133
R8343 VDD.n631 VDD.n630 1.133
R8344 VDD.n633 VDD.n632 1.133
R8345 VDD.n635 VDD.n634 1.133
R8346 VDD.n637 VDD.n636 1.133
R8347 VDD.n639 VDD.n638 1.133
R8348 VDD.n641 VDD.n640 1.133
R8349 VDD.n643 VDD.n642 1.133
R8350 VDD.n645 VDD.n644 1.133
R8351 VDD.n649 VDD.n648 1.133
R8352 VDD.n651 VDD.n650 1.133
R8353 VDD.n653 VDD.n652 1.133
R8354 VDD.n655 VDD.n654 1.133
R8355 VDD.n657 VDD.n656 1.133
R8356 VDD.n659 VDD.n658 1.133
R8357 VDD.n666 VDD.n665 1.133
R8358 VDD.n664 VDD.n663 1.133
R8359 VDD.n592 VDD.n591 1.133
R8360 VDD.n594 VDD.n593 1.133
R8361 VDD.n740 VDD.n738 1.133
R8362 VDD.n812 VDD.n810 1.133
R8363 VDD.n884 VDD.n882 1.133
R8364 VDD.n956 VDD.n954 1.133
R8365 VDD.n1028 VDD.n1026 1.133
R8366 VDD.n1100 VDD.n1098 1.133
R8367 VDD.n1172 VDD.n1170 1.133
R8368 VDD.n1244 VDD.n1242 1.133
R8369 VDD.n1316 VDD.n1314 1.133
R8370 VDD.n1388 VDD.n1386 1.133
R8371 VDD.n1460 VDD.n1458 1.133
R8372 VDD.n1532 VDD.n1530 1.133
R8373 VDD.n1604 VDD.n1602 1.133
R8374 VDD.n1676 VDD.n1675 1.133
R8375 VDD.n668 VDD.n666 1.133
R8376 VDD.n596 VDD.n594 1.133
R8377 VDD.n688 VDD.n687 0.991
R8378 VDD.n760 VDD.n759 0.991
R8379 VDD.n832 VDD.n831 0.991
R8380 VDD.n904 VDD.n903 0.991
R8381 VDD.n976 VDD.n975 0.991
R8382 VDD.n1048 VDD.n1047 0.991
R8383 VDD.n1120 VDD.n1119 0.991
R8384 VDD.n1192 VDD.n1191 0.991
R8385 VDD.n1264 VDD.n1263 0.991
R8386 VDD.n1336 VDD.n1335 0.991
R8387 VDD.n1408 VDD.n1407 0.991
R8388 VDD.n1480 VDD.n1479 0.991
R8389 VDD.n1552 VDD.n1551 0.991
R8390 VDD.n1632 VDD.n1631 0.991
R8391 VDD.n548 VDD.n547 0.991
R8392 VDD.n616 VDD.n612 0.991
R8393 VDD.n735 VDD.n731 0.964
R8394 VDD.n807 VDD.n803 0.964
R8395 VDD.n879 VDD.n875 0.964
R8396 VDD.n951 VDD.n947 0.964
R8397 VDD.n1023 VDD.n1019 0.964
R8398 VDD.n1095 VDD.n1091 0.964
R8399 VDD.n1167 VDD.n1163 0.964
R8400 VDD.n1239 VDD.n1235 0.964
R8401 VDD.n1311 VDD.n1307 0.964
R8402 VDD.n1383 VDD.n1379 0.964
R8403 VDD.n1455 VDD.n1451 0.964
R8404 VDD.n1527 VDD.n1523 0.964
R8405 VDD.n1599 VDD.n1595 0.964
R8406 VDD.n1672 VDD.n1671 0.964
R8407 VDD.n591 VDD.n587 0.964
R8408 VDD.n663 VDD.n659 0.964
R8409 VDD.n1101 VDD.n1029 0.885
R8410 VDD.n1461 VDD.n1389 0.885
R8411 VDD.n1677 VDD.n1605 0.885
R8412 VDD.n813 VDD.n741 0.884
R8413 VDD.n885 VDD.n813 0.884
R8414 VDD.n1029 VDD.n957 0.884
R8415 VDD.n1173 VDD.n1101 0.884
R8416 VDD.n1245 VDD.n1173 0.884
R8417 VDD.n1317 VDD.n1245 0.884
R8418 VDD.n1605 VDD.n1533 0.884
R8419 VDD.n741 VDD.n669 0.882
R8420 VDD.n957 VDD.n885 0.882
R8421 VDD.n1389 VDD.n1317 0.882
R8422 VDD.n1533 VDD.n1461 0.881
R8423 VDD.n702 VDD.n699 0.83
R8424 VDD.n774 VDD.n771 0.83
R8425 VDD.n846 VDD.n843 0.83
R8426 VDD.n918 VDD.n915 0.83
R8427 VDD.n990 VDD.n987 0.83
R8428 VDD.n1062 VDD.n1059 0.83
R8429 VDD.n1134 VDD.n1131 0.83
R8430 VDD.n1206 VDD.n1203 0.83
R8431 VDD.n1278 VDD.n1275 0.83
R8432 VDD.n1350 VDD.n1347 0.83
R8433 VDD.n1422 VDD.n1419 0.83
R8434 VDD.n1494 VDD.n1491 0.83
R8435 VDD.n1566 VDD.n1563 0.83
R8436 VDD.n1644 VDD.n1643 0.83
R8437 VDD.n560 VDD.n559 0.83
R8438 VDD.n630 VDD.n627 0.83
R8439 VDD.n720 VDD.n717 0.821
R8440 VDD.n792 VDD.n789 0.821
R8441 VDD.n864 VDD.n861 0.821
R8442 VDD.n936 VDD.n933 0.821
R8443 VDD.n1008 VDD.n1005 0.821
R8444 VDD.n1080 VDD.n1077 0.821
R8445 VDD.n1152 VDD.n1149 0.821
R8446 VDD.n1224 VDD.n1221 0.821
R8447 VDD.n1296 VDD.n1293 0.821
R8448 VDD.n1368 VDD.n1365 0.821
R8449 VDD.n1440 VDD.n1437 0.821
R8450 VDD.n1512 VDD.n1509 0.821
R8451 VDD.n1584 VDD.n1581 0.821
R8452 VDD.n1660 VDD.n1659 0.821
R8453 VDD.n576 VDD.n575 0.821
R8454 VDD.n648 VDD.n645 0.821
R8455 VDD.n1677 VDD.n1676 0.677
R8456 VDD.n741 VDD.n740 0.677
R8457 VDD.n813 VDD.n812 0.677
R8458 VDD.n885 VDD.n884 0.677
R8459 VDD.n1029 VDD.n1028 0.677
R8460 VDD.n1101 VDD.n1100 0.677
R8461 VDD.n1173 VDD.n1172 0.677
R8462 VDD.n1245 VDD.n1244 0.677
R8463 VDD.n1317 VDD.n1316 0.677
R8464 VDD.n1389 VDD.n1388 0.677
R8465 VDD.n1461 VDD.n1460 0.677
R8466 VDD.n1533 VDD.n1532 0.677
R8467 VDD.n1605 VDD.n1604 0.677
R8468 VDD.n669 VDD.n668 0.677
R8469 VDD.n957 VDD.n956 0.668
R8470 VDD.n690 VDD.n689 0.464
R8471 VDD.n692 VDD.n691 0.464
R8472 VDD.n694 VDD.n693 0.464
R8473 VDD.n696 VDD.n695 0.464
R8474 VDD.n698 VDD.n697 0.464
R8475 VDD.n704 VDD.n703 0.464
R8476 VDD.n706 VDD.n705 0.464
R8477 VDD.n708 VDD.n707 0.464
R8478 VDD.n710 VDD.n709 0.464
R8479 VDD.n712 VDD.n711 0.464
R8480 VDD.n714 VDD.n713 0.464
R8481 VDD.n716 VDD.n715 0.464
R8482 VDD.n722 VDD.n721 0.464
R8483 VDD.n724 VDD.n723 0.464
R8484 VDD.n726 VDD.n725 0.464
R8485 VDD.n728 VDD.n727 0.464
R8486 VDD.n730 VDD.n729 0.464
R8487 VDD.n737 VDD.n736 0.464
R8488 VDD.n686 VDD.n685 0.464
R8489 VDD.n762 VDD.n761 0.464
R8490 VDD.n764 VDD.n763 0.464
R8491 VDD.n766 VDD.n765 0.464
R8492 VDD.n768 VDD.n767 0.464
R8493 VDD.n770 VDD.n769 0.464
R8494 VDD.n776 VDD.n775 0.464
R8495 VDD.n778 VDD.n777 0.464
R8496 VDD.n780 VDD.n779 0.464
R8497 VDD.n782 VDD.n781 0.464
R8498 VDD.n784 VDD.n783 0.464
R8499 VDD.n786 VDD.n785 0.464
R8500 VDD.n788 VDD.n787 0.464
R8501 VDD.n794 VDD.n793 0.464
R8502 VDD.n796 VDD.n795 0.464
R8503 VDD.n798 VDD.n797 0.464
R8504 VDD.n800 VDD.n799 0.464
R8505 VDD.n802 VDD.n801 0.464
R8506 VDD.n809 VDD.n808 0.464
R8507 VDD.n758 VDD.n757 0.464
R8508 VDD.n834 VDD.n833 0.464
R8509 VDD.n836 VDD.n835 0.464
R8510 VDD.n838 VDD.n837 0.464
R8511 VDD.n840 VDD.n839 0.464
R8512 VDD.n842 VDD.n841 0.464
R8513 VDD.n848 VDD.n847 0.464
R8514 VDD.n850 VDD.n849 0.464
R8515 VDD.n852 VDD.n851 0.464
R8516 VDD.n854 VDD.n853 0.464
R8517 VDD.n856 VDD.n855 0.464
R8518 VDD.n858 VDD.n857 0.464
R8519 VDD.n860 VDD.n859 0.464
R8520 VDD.n866 VDD.n865 0.464
R8521 VDD.n868 VDD.n867 0.464
R8522 VDD.n870 VDD.n869 0.464
R8523 VDD.n872 VDD.n871 0.464
R8524 VDD.n874 VDD.n873 0.464
R8525 VDD.n881 VDD.n880 0.464
R8526 VDD.n830 VDD.n829 0.464
R8527 VDD.n906 VDD.n905 0.464
R8528 VDD.n908 VDD.n907 0.464
R8529 VDD.n910 VDD.n909 0.464
R8530 VDD.n912 VDD.n911 0.464
R8531 VDD.n914 VDD.n913 0.464
R8532 VDD.n920 VDD.n919 0.464
R8533 VDD.n922 VDD.n921 0.464
R8534 VDD.n924 VDD.n923 0.464
R8535 VDD.n926 VDD.n925 0.464
R8536 VDD.n928 VDD.n927 0.464
R8537 VDD.n930 VDD.n929 0.464
R8538 VDD.n932 VDD.n931 0.464
R8539 VDD.n938 VDD.n937 0.464
R8540 VDD.n940 VDD.n939 0.464
R8541 VDD.n942 VDD.n941 0.464
R8542 VDD.n944 VDD.n943 0.464
R8543 VDD.n946 VDD.n945 0.464
R8544 VDD.n953 VDD.n952 0.464
R8545 VDD.n902 VDD.n901 0.464
R8546 VDD.n978 VDD.n977 0.464
R8547 VDD.n980 VDD.n979 0.464
R8548 VDD.n982 VDD.n981 0.464
R8549 VDD.n984 VDD.n983 0.464
R8550 VDD.n986 VDD.n985 0.464
R8551 VDD.n992 VDD.n991 0.464
R8552 VDD.n994 VDD.n993 0.464
R8553 VDD.n996 VDD.n995 0.464
R8554 VDD.n998 VDD.n997 0.464
R8555 VDD.n1000 VDD.n999 0.464
R8556 VDD.n1002 VDD.n1001 0.464
R8557 VDD.n1004 VDD.n1003 0.464
R8558 VDD.n1010 VDD.n1009 0.464
R8559 VDD.n1012 VDD.n1011 0.464
R8560 VDD.n1014 VDD.n1013 0.464
R8561 VDD.n1016 VDD.n1015 0.464
R8562 VDD.n1018 VDD.n1017 0.464
R8563 VDD.n1025 VDD.n1024 0.464
R8564 VDD.n974 VDD.n973 0.464
R8565 VDD.n1050 VDD.n1049 0.464
R8566 VDD.n1052 VDD.n1051 0.464
R8567 VDD.n1054 VDD.n1053 0.464
R8568 VDD.n1056 VDD.n1055 0.464
R8569 VDD.n1058 VDD.n1057 0.464
R8570 VDD.n1064 VDD.n1063 0.464
R8571 VDD.n1066 VDD.n1065 0.464
R8572 VDD.n1068 VDD.n1067 0.464
R8573 VDD.n1070 VDD.n1069 0.464
R8574 VDD.n1072 VDD.n1071 0.464
R8575 VDD.n1074 VDD.n1073 0.464
R8576 VDD.n1076 VDD.n1075 0.464
R8577 VDD.n1082 VDD.n1081 0.464
R8578 VDD.n1084 VDD.n1083 0.464
R8579 VDD.n1086 VDD.n1085 0.464
R8580 VDD.n1088 VDD.n1087 0.464
R8581 VDD.n1090 VDD.n1089 0.464
R8582 VDD.n1097 VDD.n1096 0.464
R8583 VDD.n1046 VDD.n1045 0.464
R8584 VDD.n1122 VDD.n1121 0.464
R8585 VDD.n1124 VDD.n1123 0.464
R8586 VDD.n1126 VDD.n1125 0.464
R8587 VDD.n1128 VDD.n1127 0.464
R8588 VDD.n1130 VDD.n1129 0.464
R8589 VDD.n1136 VDD.n1135 0.464
R8590 VDD.n1138 VDD.n1137 0.464
R8591 VDD.n1140 VDD.n1139 0.464
R8592 VDD.n1142 VDD.n1141 0.464
R8593 VDD.n1144 VDD.n1143 0.464
R8594 VDD.n1146 VDD.n1145 0.464
R8595 VDD.n1148 VDD.n1147 0.464
R8596 VDD.n1154 VDD.n1153 0.464
R8597 VDD.n1156 VDD.n1155 0.464
R8598 VDD.n1158 VDD.n1157 0.464
R8599 VDD.n1160 VDD.n1159 0.464
R8600 VDD.n1162 VDD.n1161 0.464
R8601 VDD.n1169 VDD.n1168 0.464
R8602 VDD.n1118 VDD.n1117 0.464
R8603 VDD.n1194 VDD.n1193 0.464
R8604 VDD.n1196 VDD.n1195 0.464
R8605 VDD.n1198 VDD.n1197 0.464
R8606 VDD.n1200 VDD.n1199 0.464
R8607 VDD.n1202 VDD.n1201 0.464
R8608 VDD.n1208 VDD.n1207 0.464
R8609 VDD.n1210 VDD.n1209 0.464
R8610 VDD.n1212 VDD.n1211 0.464
R8611 VDD.n1214 VDD.n1213 0.464
R8612 VDD.n1216 VDD.n1215 0.464
R8613 VDD.n1218 VDD.n1217 0.464
R8614 VDD.n1220 VDD.n1219 0.464
R8615 VDD.n1226 VDD.n1225 0.464
R8616 VDD.n1228 VDD.n1227 0.464
R8617 VDD.n1230 VDD.n1229 0.464
R8618 VDD.n1232 VDD.n1231 0.464
R8619 VDD.n1234 VDD.n1233 0.464
R8620 VDD.n1241 VDD.n1240 0.464
R8621 VDD.n1190 VDD.n1189 0.464
R8622 VDD.n1266 VDD.n1265 0.464
R8623 VDD.n1268 VDD.n1267 0.464
R8624 VDD.n1270 VDD.n1269 0.464
R8625 VDD.n1272 VDD.n1271 0.464
R8626 VDD.n1274 VDD.n1273 0.464
R8627 VDD.n1280 VDD.n1279 0.464
R8628 VDD.n1282 VDD.n1281 0.464
R8629 VDD.n1284 VDD.n1283 0.464
R8630 VDD.n1286 VDD.n1285 0.464
R8631 VDD.n1288 VDD.n1287 0.464
R8632 VDD.n1290 VDD.n1289 0.464
R8633 VDD.n1292 VDD.n1291 0.464
R8634 VDD.n1298 VDD.n1297 0.464
R8635 VDD.n1300 VDD.n1299 0.464
R8636 VDD.n1302 VDD.n1301 0.464
R8637 VDD.n1304 VDD.n1303 0.464
R8638 VDD.n1306 VDD.n1305 0.464
R8639 VDD.n1313 VDD.n1312 0.464
R8640 VDD.n1262 VDD.n1261 0.464
R8641 VDD.n1338 VDD.n1337 0.464
R8642 VDD.n1340 VDD.n1339 0.464
R8643 VDD.n1342 VDD.n1341 0.464
R8644 VDD.n1344 VDD.n1343 0.464
R8645 VDD.n1346 VDD.n1345 0.464
R8646 VDD.n1352 VDD.n1351 0.464
R8647 VDD.n1354 VDD.n1353 0.464
R8648 VDD.n1356 VDD.n1355 0.464
R8649 VDD.n1358 VDD.n1357 0.464
R8650 VDD.n1360 VDD.n1359 0.464
R8651 VDD.n1362 VDD.n1361 0.464
R8652 VDD.n1364 VDD.n1363 0.464
R8653 VDD.n1370 VDD.n1369 0.464
R8654 VDD.n1372 VDD.n1371 0.464
R8655 VDD.n1374 VDD.n1373 0.464
R8656 VDD.n1376 VDD.n1375 0.464
R8657 VDD.n1378 VDD.n1377 0.464
R8658 VDD.n1385 VDD.n1384 0.464
R8659 VDD.n1334 VDD.n1333 0.464
R8660 VDD.n1410 VDD.n1409 0.464
R8661 VDD.n1412 VDD.n1411 0.464
R8662 VDD.n1414 VDD.n1413 0.464
R8663 VDD.n1416 VDD.n1415 0.464
R8664 VDD.n1418 VDD.n1417 0.464
R8665 VDD.n1424 VDD.n1423 0.464
R8666 VDD.n1426 VDD.n1425 0.464
R8667 VDD.n1428 VDD.n1427 0.464
R8668 VDD.n1430 VDD.n1429 0.464
R8669 VDD.n1432 VDD.n1431 0.464
R8670 VDD.n1434 VDD.n1433 0.464
R8671 VDD.n1436 VDD.n1435 0.464
R8672 VDD.n1442 VDD.n1441 0.464
R8673 VDD.n1444 VDD.n1443 0.464
R8674 VDD.n1446 VDD.n1445 0.464
R8675 VDD.n1448 VDD.n1447 0.464
R8676 VDD.n1450 VDD.n1449 0.464
R8677 VDD.n1457 VDD.n1456 0.464
R8678 VDD.n1406 VDD.n1405 0.464
R8679 VDD.n1482 VDD.n1481 0.464
R8680 VDD.n1484 VDD.n1483 0.464
R8681 VDD.n1486 VDD.n1485 0.464
R8682 VDD.n1488 VDD.n1487 0.464
R8683 VDD.n1490 VDD.n1489 0.464
R8684 VDD.n1496 VDD.n1495 0.464
R8685 VDD.n1498 VDD.n1497 0.464
R8686 VDD.n1500 VDD.n1499 0.464
R8687 VDD.n1502 VDD.n1501 0.464
R8688 VDD.n1504 VDD.n1503 0.464
R8689 VDD.n1506 VDD.n1505 0.464
R8690 VDD.n1508 VDD.n1507 0.464
R8691 VDD.n1514 VDD.n1513 0.464
R8692 VDD.n1516 VDD.n1515 0.464
R8693 VDD.n1518 VDD.n1517 0.464
R8694 VDD.n1520 VDD.n1519 0.464
R8695 VDD.n1522 VDD.n1521 0.464
R8696 VDD.n1529 VDD.n1528 0.464
R8697 VDD.n1478 VDD.n1477 0.464
R8698 VDD.n1554 VDD.n1553 0.464
R8699 VDD.n1556 VDD.n1555 0.464
R8700 VDD.n1558 VDD.n1557 0.464
R8701 VDD.n1560 VDD.n1559 0.464
R8702 VDD.n1562 VDD.n1561 0.464
R8703 VDD.n1568 VDD.n1567 0.464
R8704 VDD.n1570 VDD.n1569 0.464
R8705 VDD.n1572 VDD.n1571 0.464
R8706 VDD.n1574 VDD.n1573 0.464
R8707 VDD.n1576 VDD.n1575 0.464
R8708 VDD.n1578 VDD.n1577 0.464
R8709 VDD.n1580 VDD.n1579 0.464
R8710 VDD.n1586 VDD.n1585 0.464
R8711 VDD.n1588 VDD.n1587 0.464
R8712 VDD.n1590 VDD.n1589 0.464
R8713 VDD.n1592 VDD.n1591 0.464
R8714 VDD.n1594 VDD.n1593 0.464
R8715 VDD.n1601 VDD.n1600 0.464
R8716 VDD.n1550 VDD.n1549 0.464
R8717 VDD.n1674 VDD.n1673 0.464
R8718 VDD.n1670 VDD.n1669 0.464
R8719 VDD.n1668 VDD.n1667 0.464
R8720 VDD.n1666 VDD.n1665 0.464
R8721 VDD.n1664 VDD.n1663 0.464
R8722 VDD.n1662 VDD.n1661 0.464
R8723 VDD.n1658 VDD.n1657 0.464
R8724 VDD.n1656 VDD.n1655 0.464
R8725 VDD.n1654 VDD.n1653 0.464
R8726 VDD.n1652 VDD.n1651 0.464
R8727 VDD.n1650 VDD.n1649 0.464
R8728 VDD.n1648 VDD.n1647 0.464
R8729 VDD.n1646 VDD.n1645 0.464
R8730 VDD.n1642 VDD.n1641 0.464
R8731 VDD.n1640 VDD.n1639 0.464
R8732 VDD.n1638 VDD.n1637 0.464
R8733 VDD.n1636 VDD.n1635 0.464
R8734 VDD.n1634 VDD.n1633 0.464
R8735 VDD.n1630 VDD.n1629 0.464
R8736 VDD.n586 VDD.n585 0.464
R8737 VDD.n584 VDD.n583 0.464
R8738 VDD.n582 VDD.n581 0.464
R8739 VDD.n580 VDD.n579 0.464
R8740 VDD.n578 VDD.n577 0.464
R8741 VDD.n574 VDD.n573 0.464
R8742 VDD.n572 VDD.n571 0.464
R8743 VDD.n570 VDD.n569 0.464
R8744 VDD.n568 VDD.n567 0.464
R8745 VDD.n566 VDD.n565 0.464
R8746 VDD.n564 VDD.n563 0.464
R8747 VDD.n562 VDD.n561 0.464
R8748 VDD.n558 VDD.n557 0.464
R8749 VDD.n556 VDD.n555 0.464
R8750 VDD.n554 VDD.n553 0.464
R8751 VDD.n552 VDD.n551 0.464
R8752 VDD.n550 VDD.n549 0.464
R8753 VDD.n546 VDD.n545 0.464
R8754 VDD.n611 VDD.n610 0.464
R8755 VDD.n618 VDD.n617 0.464
R8756 VDD.n620 VDD.n619 0.464
R8757 VDD.n622 VDD.n621 0.464
R8758 VDD.n624 VDD.n623 0.464
R8759 VDD.n626 VDD.n625 0.464
R8760 VDD.n632 VDD.n631 0.464
R8761 VDD.n634 VDD.n633 0.464
R8762 VDD.n636 VDD.n635 0.464
R8763 VDD.n638 VDD.n637 0.464
R8764 VDD.n640 VDD.n639 0.464
R8765 VDD.n642 VDD.n641 0.464
R8766 VDD.n644 VDD.n643 0.464
R8767 VDD.n650 VDD.n649 0.464
R8768 VDD.n652 VDD.n651 0.464
R8769 VDD.n654 VDD.n653 0.464
R8770 VDD.n656 VDD.n655 0.464
R8771 VDD.n658 VDD.n657 0.464
R8772 VDD.n665 VDD.n664 0.464
R8773 VDD.n593 VDD.n592 0.464
R8774 VDD VDD.n1678 0.367
R8775 VDD.n27 VDD.n25 0.042
R8776 VDD.n12 VDD.n10 0.042
R8777 VDD.n19 VDD.n18 0.042
R8778 VDD.n18 VDD.n17 0.042
R8779 VDD.n31 VDD.n30 0.042
R8780 VDD.n30 VDD.n29 0.042
R8781 VDD.n59 VDD.n57 0.042
R8782 VDD.n44 VDD.n42 0.042
R8783 VDD.n51 VDD.n50 0.042
R8784 VDD.n50 VDD.n49 0.042
R8785 VDD.n63 VDD.n62 0.042
R8786 VDD.n62 VDD.n61 0.042
R8787 VDD.n91 VDD.n89 0.042
R8788 VDD.n76 VDD.n74 0.042
R8789 VDD.n83 VDD.n82 0.042
R8790 VDD.n82 VDD.n81 0.042
R8791 VDD.n95 VDD.n94 0.042
R8792 VDD.n94 VDD.n93 0.042
R8793 VDD.n123 VDD.n121 0.042
R8794 VDD.n108 VDD.n106 0.042
R8795 VDD.n115 VDD.n114 0.042
R8796 VDD.n114 VDD.n113 0.042
R8797 VDD.n127 VDD.n126 0.042
R8798 VDD.n126 VDD.n125 0.042
R8799 VDD.n155 VDD.n153 0.042
R8800 VDD.n140 VDD.n138 0.042
R8801 VDD.n147 VDD.n146 0.042
R8802 VDD.n146 VDD.n145 0.042
R8803 VDD.n159 VDD.n158 0.042
R8804 VDD.n158 VDD.n157 0.042
R8805 VDD.n187 VDD.n185 0.042
R8806 VDD.n172 VDD.n170 0.042
R8807 VDD.n179 VDD.n178 0.042
R8808 VDD.n178 VDD.n177 0.042
R8809 VDD.n191 VDD.n190 0.042
R8810 VDD.n190 VDD.n189 0.042
R8811 VDD.n219 VDD.n217 0.042
R8812 VDD.n204 VDD.n202 0.042
R8813 VDD.n211 VDD.n210 0.042
R8814 VDD.n210 VDD.n209 0.042
R8815 VDD.n223 VDD.n222 0.042
R8816 VDD.n222 VDD.n221 0.042
R8817 VDD.n251 VDD.n249 0.042
R8818 VDD.n236 VDD.n234 0.042
R8819 VDD.n243 VDD.n242 0.042
R8820 VDD.n242 VDD.n241 0.042
R8821 VDD.n255 VDD.n254 0.042
R8822 VDD.n254 VDD.n253 0.042
R8823 VDD.n283 VDD.n281 0.042
R8824 VDD.n268 VDD.n266 0.042
R8825 VDD.n275 VDD.n274 0.042
R8826 VDD.n274 VDD.n273 0.042
R8827 VDD.n287 VDD.n286 0.042
R8828 VDD.n286 VDD.n285 0.042
R8829 VDD.n315 VDD.n313 0.042
R8830 VDD.n300 VDD.n298 0.042
R8831 VDD.n307 VDD.n306 0.042
R8832 VDD.n306 VDD.n305 0.042
R8833 VDD.n319 VDD.n318 0.042
R8834 VDD.n318 VDD.n317 0.042
R8835 VDD.n347 VDD.n345 0.042
R8836 VDD.n332 VDD.n330 0.042
R8837 VDD.n339 VDD.n338 0.042
R8838 VDD.n338 VDD.n337 0.042
R8839 VDD.n351 VDD.n350 0.042
R8840 VDD.n350 VDD.n349 0.042
R8841 VDD.n379 VDD.n377 0.042
R8842 VDD.n364 VDD.n362 0.042
R8843 VDD.n371 VDD.n370 0.042
R8844 VDD.n370 VDD.n369 0.042
R8845 VDD.n383 VDD.n382 0.042
R8846 VDD.n382 VDD.n381 0.042
R8847 VDD.n411 VDD.n409 0.042
R8848 VDD.n396 VDD.n394 0.042
R8849 VDD.n403 VDD.n402 0.042
R8850 VDD.n402 VDD.n401 0.042
R8851 VDD.n415 VDD.n414 0.042
R8852 VDD.n414 VDD.n413 0.042
R8853 VDD.n443 VDD.n441 0.042
R8854 VDD.n428 VDD.n426 0.042
R8855 VDD.n435 VDD.n434 0.042
R8856 VDD.n434 VDD.n433 0.042
R8857 VDD.n447 VDD.n446 0.042
R8858 VDD.n446 VDD.n445 0.042
R8859 VDD.n475 VDD.n473 0.042
R8860 VDD.n460 VDD.n458 0.042
R8861 VDD.n467 VDD.n466 0.042
R8862 VDD.n466 VDD.n465 0.042
R8863 VDD.n479 VDD.n478 0.042
R8864 VDD.n478 VDD.n477 0.042
R8865 VDD.n507 VDD.n505 0.042
R8866 VDD.n492 VDD.n490 0.042
R8867 VDD.n499 VDD.n498 0.042
R8868 VDD.n498 VDD.n497 0.042
R8869 VDD.n511 VDD.n510 0.042
R8870 VDD.n510 VDD.n509 0.042
R8871 VDD.n599 VDD.n597 0.042
R8872 VDD.n675 VDD.n673 0.042
R8873 VDD.n683 VDD.n682 0.042
R8874 VDD.n682 VDD.n681 0.042
R8875 VDD.n747 VDD.n745 0.042
R8876 VDD.n755 VDD.n754 0.042
R8877 VDD.n754 VDD.n753 0.042
R8878 VDD.n819 VDD.n817 0.042
R8879 VDD.n827 VDD.n826 0.042
R8880 VDD.n826 VDD.n825 0.042
R8881 VDD.n891 VDD.n889 0.042
R8882 VDD.n899 VDD.n898 0.042
R8883 VDD.n898 VDD.n897 0.042
R8884 VDD.n963 VDD.n961 0.042
R8885 VDD.n971 VDD.n970 0.042
R8886 VDD.n970 VDD.n969 0.042
R8887 VDD.n1035 VDD.n1033 0.042
R8888 VDD.n1043 VDD.n1042 0.042
R8889 VDD.n1042 VDD.n1041 0.042
R8890 VDD.n1107 VDD.n1105 0.042
R8891 VDD.n1115 VDD.n1114 0.042
R8892 VDD.n1114 VDD.n1113 0.042
R8893 VDD.n1179 VDD.n1177 0.042
R8894 VDD.n1187 VDD.n1186 0.042
R8895 VDD.n1186 VDD.n1185 0.042
R8896 VDD.n1251 VDD.n1249 0.042
R8897 VDD.n1259 VDD.n1258 0.042
R8898 VDD.n1258 VDD.n1257 0.042
R8899 VDD.n1323 VDD.n1321 0.042
R8900 VDD.n1331 VDD.n1330 0.042
R8901 VDD.n1330 VDD.n1329 0.042
R8902 VDD.n1395 VDD.n1393 0.042
R8903 VDD.n1403 VDD.n1402 0.042
R8904 VDD.n1402 VDD.n1401 0.042
R8905 VDD.n1467 VDD.n1465 0.042
R8906 VDD.n1475 VDD.n1474 0.042
R8907 VDD.n1474 VDD.n1473 0.042
R8908 VDD.n1539 VDD.n1537 0.042
R8909 VDD.n1547 VDD.n1546 0.042
R8910 VDD.n1546 VDD.n1545 0.042
R8911 VDD.n1619 VDD.n1617 0.042
R8912 VDD.n1627 VDD.n1626 0.042
R8913 VDD.n1626 VDD.n1625 0.042
R8914 VDD.n536 VDD.n534 0.042
R8915 VDD.n543 VDD.n542 0.042
R8916 VDD.n542 VDD.n541 0.042
R8917 VDD.n608 VDD.n607 0.042
R8918 VDD.n607 VDD.n606 0.042
R8919 VDD.n21 VDD.n20 0.039
R8920 VDD.n53 VDD.n52 0.039
R8921 VDD.n85 VDD.n84 0.039
R8922 VDD.n117 VDD.n116 0.039
R8923 VDD.n149 VDD.n148 0.039
R8924 VDD.n181 VDD.n180 0.039
R8925 VDD.n213 VDD.n212 0.039
R8926 VDD.n245 VDD.n244 0.039
R8927 VDD.n277 VDD.n276 0.039
R8928 VDD.n309 VDD.n308 0.039
R8929 VDD.n341 VDD.n340 0.039
R8930 VDD.n373 VDD.n372 0.039
R8931 VDD.n405 VDD.n404 0.039
R8932 VDD.n437 VDD.n436 0.039
R8933 VDD.n469 VDD.n468 0.039
R8934 VDD.n501 VDD.n500 0.039
R8935 VDD.n16 VDD.n15 0.023
R8936 VDD.n28 VDD.n21 0.023
R8937 VDD.n48 VDD.n47 0.023
R8938 VDD.n60 VDD.n53 0.023
R8939 VDD.n80 VDD.n79 0.023
R8940 VDD.n92 VDD.n85 0.023
R8941 VDD.n112 VDD.n111 0.023
R8942 VDD.n124 VDD.n117 0.023
R8943 VDD.n144 VDD.n143 0.023
R8944 VDD.n156 VDD.n149 0.023
R8945 VDD.n176 VDD.n175 0.023
R8946 VDD.n188 VDD.n181 0.023
R8947 VDD.n208 VDD.n207 0.023
R8948 VDD.n220 VDD.n213 0.023
R8949 VDD.n240 VDD.n239 0.023
R8950 VDD.n252 VDD.n245 0.023
R8951 VDD.n272 VDD.n271 0.023
R8952 VDD.n284 VDD.n277 0.023
R8953 VDD.n304 VDD.n303 0.023
R8954 VDD.n316 VDD.n309 0.023
R8955 VDD.n336 VDD.n335 0.023
R8956 VDD.n348 VDD.n341 0.023
R8957 VDD.n368 VDD.n367 0.023
R8958 VDD.n380 VDD.n373 0.023
R8959 VDD.n400 VDD.n399 0.023
R8960 VDD.n412 VDD.n405 0.023
R8961 VDD.n432 VDD.n431 0.023
R8962 VDD.n444 VDD.n437 0.023
R8963 VDD.n464 VDD.n463 0.023
R8964 VDD.n476 VDD.n469 0.023
R8965 VDD.n496 VDD.n495 0.023
R8966 VDD.n508 VDD.n501 0.023
R8967 VDD.n7 VDD.n6 0.021
R8968 VDD.n27 VDD.n24 0.021
R8969 VDD.n4 VDD.n2 0.021
R8970 VDD.n41 VDD.n39 0.021
R8971 VDD.n59 VDD.n56 0.021
R8972 VDD.n34 VDD.n33 0.021
R8973 VDD.n71 VDD.n70 0.021
R8974 VDD.n91 VDD.n88 0.021
R8975 VDD.n68 VDD.n66 0.021
R8976 VDD.n103 VDD.n102 0.021
R8977 VDD.n123 VDD.n120 0.021
R8978 VDD.n98 VDD.n97 0.021
R8979 VDD.n135 VDD.n134 0.021
R8980 VDD.n155 VDD.n152 0.021
R8981 VDD.n130 VDD.n129 0.021
R8982 VDD.n169 VDD.n167 0.021
R8983 VDD.n187 VDD.n184 0.021
R8984 VDD.n164 VDD.n162 0.021
R8985 VDD.n199 VDD.n198 0.021
R8986 VDD.n219 VDD.n216 0.021
R8987 VDD.n194 VDD.n193 0.021
R8988 VDD.n231 VDD.n230 0.021
R8989 VDD.n251 VDD.n248 0.021
R8990 VDD.n226 VDD.n225 0.021
R8991 VDD.n265 VDD.n263 0.021
R8992 VDD.n283 VDD.n280 0.021
R8993 VDD.n258 VDD.n257 0.021
R8994 VDD.n295 VDD.n294 0.021
R8995 VDD.n315 VDD.n312 0.021
R8996 VDD.n290 VDD.n289 0.021
R8997 VDD.n329 VDD.n327 0.021
R8998 VDD.n347 VDD.n344 0.021
R8999 VDD.n322 VDD.n321 0.021
R9000 VDD.n359 VDD.n358 0.021
R9001 VDD.n379 VDD.n376 0.021
R9002 VDD.n356 VDD.n354 0.021
R9003 VDD.n393 VDD.n391 0.021
R9004 VDD.n411 VDD.n408 0.021
R9005 VDD.n388 VDD.n386 0.021
R9006 VDD.n423 VDD.n422 0.021
R9007 VDD.n443 VDD.n440 0.021
R9008 VDD.n420 VDD.n418 0.021
R9009 VDD.n457 VDD.n455 0.021
R9010 VDD.n475 VDD.n472 0.021
R9011 VDD.n450 VDD.n449 0.021
R9012 VDD.n487 VDD.n486 0.021
R9013 VDD.n507 VDD.n504 0.021
R9014 VDD.n484 VDD.n482 0.021
R9015 VDD.n14 VDD.n12 0.015
R9016 VDD.n46 VDD.n44 0.015
R9017 VDD.n78 VDD.n76 0.015
R9018 VDD.n110 VDD.n108 0.015
R9019 VDD.n142 VDD.n140 0.015
R9020 VDD.n174 VDD.n172 0.015
R9021 VDD.n206 VDD.n204 0.015
R9022 VDD.n238 VDD.n236 0.015
R9023 VDD.n270 VDD.n268 0.015
R9024 VDD.n302 VDD.n300 0.015
R9025 VDD.n334 VDD.n332 0.015
R9026 VDD.n366 VDD.n364 0.015
R9027 VDD.n398 VDD.n396 0.015
R9028 VDD.n430 VDD.n428 0.015
R9029 VDD.n462 VDD.n460 0.015
R9030 VDD.n494 VDD.n492 0.015
R9031 VDD.n676 VDD.n675 0.015
R9032 VDD.n748 VDD.n747 0.015
R9033 VDD.n820 VDD.n819 0.015
R9034 VDD.n892 VDD.n891 0.015
R9035 VDD.n964 VDD.n963 0.015
R9036 VDD.n1036 VDD.n1035 0.015
R9037 VDD.n1108 VDD.n1107 0.015
R9038 VDD.n1180 VDD.n1179 0.015
R9039 VDD.n1252 VDD.n1251 0.015
R9040 VDD.n1324 VDD.n1323 0.015
R9041 VDD.n1396 VDD.n1395 0.015
R9042 VDD.n1468 VDD.n1467 0.015
R9043 VDD.n1540 VDD.n1539 0.015
R9044 VDD.n1620 VDD.n1619 0.015
R9045 VDD.n537 VDD.n536 0.015
R9046 VDD.n600 VDD.n599 0.015
R9047 SA_OUT[5].n0 SA_OUT[5].t4 661.027
R9048 SA_OUT[5].n0 SA_OUT[5].t3 392.255
R9049 SA_OUT[5].n1 SA_OUT[5].t1 223.716
R9050 SA_OUT[5].n2 SA_OUT[5].t0 153.977
R9051 SA_OUT[5].n1 SA_OUT[5].n0 143.764
R9052 SA_OUT[5].n2 SA_OUT[5].t2 59.86
R9053 SA_OUT[5] SA_OUT[5].n2 17.544
R9054 SA_OUT[5].n2 SA_OUT[5].n1 4.517
R9055 a_8340_n812.t0 a_8340_n812.t1 242.857
R9056 a_8340_n953.t35 a_8340_n953.n46 176.385
R9057 a_8340_n953.n22 a_8340_n953.t14 67.378
R9058 a_8340_n953.n0 a_8340_n953.t19 66.92
R9059 a_8340_n953.n1 a_8340_n953.t11 66.92
R9060 a_8340_n953.n2 a_8340_n953.t18 66.92
R9061 a_8340_n953.n3 a_8340_n953.t9 66.92
R9062 a_8340_n953.n4 a_8340_n953.t5 66.92
R9063 a_8340_n953.n5 a_8340_n953.t48 66.92
R9064 a_8340_n953.n6 a_8340_n953.t37 66.92
R9065 a_8340_n953.n7 a_8340_n953.t41 66.92
R9066 a_8340_n953.n8 a_8340_n953.t26 66.92
R9067 a_8340_n953.n9 a_8340_n953.t1 66.92
R9068 a_8340_n953.n10 a_8340_n953.t22 66.92
R9069 a_8340_n953.n11 a_8340_n953.t31 66.92
R9070 a_8340_n953.n12 a_8340_n953.t28 66.92
R9071 a_8340_n953.n13 a_8340_n953.t43 66.92
R9072 a_8340_n953.n14 a_8340_n953.t47 66.92
R9073 a_8340_n953.n15 a_8340_n953.t45 66.92
R9074 a_8340_n953.n16 a_8340_n953.t39 66.92
R9075 a_8340_n953.n17 a_8340_n953.t0 66.92
R9076 a_8340_n953.n18 a_8340_n953.t25 66.92
R9077 a_8340_n953.n19 a_8340_n953.t46 66.92
R9078 a_8340_n953.n20 a_8340_n953.t15 66.92
R9079 a_8340_n953.n21 a_8340_n953.t16 66.92
R9080 a_8340_n953.n22 a_8340_n953.t21 66.92
R9081 a_8340_n953.n23 a_8340_n953.t6 65.518
R9082 a_8340_n953.n45 a_8340_n953.t7 63.519
R9083 a_8340_n953.n44 a_8340_n953.t20 63.519
R9084 a_8340_n953.n43 a_8340_n953.t10 63.519
R9085 a_8340_n953.n42 a_8340_n953.t12 63.519
R9086 a_8340_n953.n41 a_8340_n953.t33 63.519
R9087 a_8340_n953.n40 a_8340_n953.t36 63.519
R9088 a_8340_n953.n39 a_8340_n953.t24 63.519
R9089 a_8340_n953.n38 a_8340_n953.t23 63.519
R9090 a_8340_n953.n37 a_8340_n953.t40 63.519
R9091 a_8340_n953.n36 a_8340_n953.t34 63.519
R9092 a_8340_n953.n35 a_8340_n953.t30 63.519
R9093 a_8340_n953.n34 a_8340_n953.t29 63.519
R9094 a_8340_n953.n33 a_8340_n953.t3 63.519
R9095 a_8340_n953.n32 a_8340_n953.t38 63.519
R9096 a_8340_n953.n31 a_8340_n953.t42 63.519
R9097 a_8340_n953.n30 a_8340_n953.t4 63.519
R9098 a_8340_n953.n29 a_8340_n953.t32 63.519
R9099 a_8340_n953.n28 a_8340_n953.t44 63.519
R9100 a_8340_n953.n27 a_8340_n953.t2 63.519
R9101 a_8340_n953.n26 a_8340_n953.t27 63.519
R9102 a_8340_n953.n25 a_8340_n953.t8 63.519
R9103 a_8340_n953.n24 a_8340_n953.t13 63.519
R9104 a_8340_n953.n23 a_8340_n953.t17 63.519
R9105 a_8340_n953.n46 a_8340_n953.n0 19.599
R9106 a_8340_n953.n46 a_8340_n953.n45 15.67
R9107 a_8340_n953.n44 a_8340_n953.n43 2.524
R9108 a_8340_n953.n24 a_8340_n953.n23 2.498
R9109 a_8340_n953.n21 a_8340_n953.n22 2.495
R9110 a_8340_n953.n1 a_8340_n953.n2 2.459
R9111 a_8340_n953.n38 a_8340_n953.n37 2.364
R9112 a_8340_n953.n30 a_8340_n953.n29 2.355
R9113 a_8340_n953.n7 a_8340_n953.n8 2.299
R9114 a_8340_n953.n15 a_8340_n953.n16 2.29
R9115 a_8340_n953.n16 a_8340_n953.n17 2.057
R9116 a_8340_n953.n8 a_8340_n953.n9 2.057
R9117 a_8340_n953.n2 a_8340_n953.n3 2.057
R9118 a_8340_n953.n0 a_8340_n953.n1 2.057
R9119 a_8340_n953.n45 a_8340_n953.n44 1.998
R9120 a_8340_n953.n43 a_8340_n953.n42 1.998
R9121 a_8340_n953.n42 a_8340_n953.n41 1.998
R9122 a_8340_n953.n41 a_8340_n953.n40 1.998
R9123 a_8340_n953.n40 a_8340_n953.n39 1.998
R9124 a_8340_n953.n39 a_8340_n953.n38 1.998
R9125 a_8340_n953.n37 a_8340_n953.n36 1.998
R9126 a_8340_n953.n36 a_8340_n953.n35 1.998
R9127 a_8340_n953.n35 a_8340_n953.n34 1.998
R9128 a_8340_n953.n34 a_8340_n953.n33 1.998
R9129 a_8340_n953.n33 a_8340_n953.n32 1.998
R9130 a_8340_n953.n32 a_8340_n953.n31 1.998
R9131 a_8340_n953.n31 a_8340_n953.n30 1.998
R9132 a_8340_n953.n29 a_8340_n953.n28 1.998
R9133 a_8340_n953.n28 a_8340_n953.n27 1.998
R9134 a_8340_n953.n27 a_8340_n953.n26 1.998
R9135 a_8340_n953.n26 a_8340_n953.n25 1.998
R9136 a_8340_n953.n25 a_8340_n953.n24 1.998
R9137 a_8340_n953.n20 a_8340_n953.n21 1.995
R9138 a_8340_n953.n19 a_8340_n953.n20 1.995
R9139 a_8340_n953.n18 a_8340_n953.n19 1.995
R9140 a_8340_n953.n17 a_8340_n953.n18 1.995
R9141 a_8340_n953.n14 a_8340_n953.n15 1.995
R9142 a_8340_n953.n13 a_8340_n953.n14 1.995
R9143 a_8340_n953.n12 a_8340_n953.n13 1.995
R9144 a_8340_n953.n11 a_8340_n953.n12 1.995
R9145 a_8340_n953.n10 a_8340_n953.n11 1.995
R9146 a_8340_n953.n9 a_8340_n953.n10 1.995
R9147 a_8340_n953.n6 a_8340_n953.n7 1.995
R9148 a_8340_n953.n5 a_8340_n953.n6 1.995
R9149 a_8340_n953.n4 a_8340_n953.n5 1.995
R9150 a_8340_n953.n3 a_8340_n953.n4 1.995
R9151 a_3247_3666.n0 a_3247_3666.t0 358.166
R9152 a_3247_3666.t4 a_3247_3666.t5 337.399
R9153 a_3247_3666.t5 a_3247_3666.t3 285.986
R9154 a_3247_3666.n0 a_3247_3666.t4 282.573
R9155 a_3247_3666.n1 a_3247_3666.t2 202.857
R9156 a_3247_3666.n1 a_3247_3666.n0 173.817
R9157 a_3247_3666.n1 a_3247_3666.t1 20.826
R9158 a_3247_3666.n2 a_3247_3666.n1 20.689
R9159 a_3617_3666.t0 a_3617_3666.t1 242.857
R9160 a_4397_1698.n0 a_4397_1698.t2 358.166
R9161 a_4397_1698.t4 a_4397_1698.t5 337.399
R9162 a_4397_1698.t5 a_4397_1698.t3 285.986
R9163 a_4397_1698.n0 a_4397_1698.t4 282.573
R9164 a_4397_1698.n1 a_4397_1698.t0 202.857
R9165 a_4397_1698.n1 a_4397_1698.n0 173.817
R9166 a_4397_1698.n1 a_4397_1698.t1 20.826
R9167 a_4397_1698.n2 a_4397_1698.n1 20.689
R9168 a_4767_1698.t0 a_4767_1698.t1 242.857
R9169 a_1427_437.n0 a_1427_437.t0 362.857
R9170 a_1427_437.t5 a_1427_437.t4 337.399
R9171 a_1427_437.t4 a_1427_437.t3 298.839
R9172 a_1427_437.n0 a_1427_437.t5 280.405
R9173 a_1427_437.n1 a_1427_437.t2 200
R9174 a_1427_437.n1 a_1427_437.n0 172.311
R9175 a_1427_437.n2 a_1427_437.n1 24
R9176 a_1427_437.n1 a_1427_437.t1 21.212
R9177 a_1440_452.t0 a_1440_452.t1 242.857
R9178 a_277_1201.n0 a_277_1201.t1 362.857
R9179 a_277_1201.t5 a_277_1201.t3 337.399
R9180 a_277_1201.t3 a_277_1201.t4 298.839
R9181 a_277_1201.n0 a_277_1201.t5 280.405
R9182 a_277_1201.n1 a_277_1201.t0 200
R9183 a_277_1201.n1 a_277_1201.n0 172.311
R9184 a_277_1201.n2 a_277_1201.n1 24
R9185 a_277_1201.n1 a_277_1201.t2 21.212
R9186 a_372_1216.n0 a_372_1216.t2 358.166
R9187 a_372_1216.t3 a_372_1216.t5 337.399
R9188 a_372_1216.t5 a_372_1216.t4 285.986
R9189 a_372_1216.n0 a_372_1216.t3 282.573
R9190 a_372_1216.n1 a_372_1216.t0 202.857
R9191 a_372_1216.n1 a_372_1216.n0 173.817
R9192 a_372_1216.n1 a_372_1216.t1 20.826
R9193 a_372_1216.n2 a_372_1216.n1 20.689
R9194 a_7827_n2234.n2 a_7827_n2234.t1 282.97
R9195 a_7827_n2234.n1 a_7827_n2234.t3 240.683
R9196 a_7827_n2234.n0 a_7827_n2234.t4 209.208
R9197 a_7827_n2234.n0 a_7827_n2234.t2 194.167
R9198 a_7827_n2234.t0 a_7827_n2234.n2 183.404
R9199 a_7827_n2234.n1 a_7827_n2234.n0 14.805
R9200 a_7827_n2234.n2 a_7827_n2234.n1 6.415
R9201 a_7950_n2132.n0 a_7950_n2132.t2 489.336
R9202 a_7950_n2132.n0 a_7950_n2132.t1 243.258
R9203 a_7950_n2132.t0 a_7950_n2132.n0 214.415
R9204 a_3247_n512.n0 a_3247_n512.t0 358.166
R9205 a_3247_n512.t5 a_3247_n512.t3 337.399
R9206 a_3247_n512.t3 a_3247_n512.t4 285.986
R9207 a_3247_n512.n0 a_3247_n512.t5 282.573
R9208 a_3247_n512.n1 a_3247_n512.t2 202.857
R9209 a_3247_n512.n1 a_3247_n512.n0 173.817
R9210 a_3247_n512.n1 a_3247_n512.t1 20.826
R9211 a_3247_n512.n2 a_3247_n512.n1 20.689
R9212 a_3152_n527.n0 a_3152_n527.t2 362.857
R9213 a_3152_n527.t3 a_3152_n527.t4 337.399
R9214 a_3152_n527.t4 a_3152_n527.t5 298.839
R9215 a_3152_n527.n0 a_3152_n527.t3 280.405
R9216 a_3152_n527.n1 a_3152_n527.t0 200
R9217 a_3152_n527.n1 a_3152_n527.n0 172.311
R9218 a_3152_n527.n2 a_3152_n527.n1 24
R9219 a_3152_n527.n1 a_3152_n527.t1 21.212
R9220 a_2002_4133.n0 a_2002_4133.t0 362.857
R9221 a_2002_4133.t3 a_2002_4133.t5 337.399
R9222 a_2002_4133.t5 a_2002_4133.t4 298.839
R9223 a_2002_4133.n0 a_2002_4133.t3 280.405
R9224 a_2002_4133.n1 a_2002_4133.t2 200
R9225 a_2002_4133.n1 a_2002_4133.n0 172.311
R9226 a_2002_4133.n2 a_2002_4133.n1 24
R9227 a_2002_4133.n1 a_2002_4133.t1 21.212
R9228 a_2097_4148.n0 a_2097_4148.t1 358.166
R9229 a_2097_4148.t5 a_2097_4148.t3 337.399
R9230 a_2097_4148.t3 a_2097_4148.t4 285.986
R9231 a_2097_4148.n0 a_2097_4148.t5 282.573
R9232 a_2097_4148.n1 a_2097_4148.t2 202.857
R9233 a_2097_4148.n1 a_2097_4148.n0 173.817
R9234 a_2097_4148.n1 a_2097_4148.t0 20.826
R9235 a_2097_4148.n2 a_2097_4148.n1 20.689
R9236 a_8327_3169.n0 a_8327_3169.t1 362.857
R9237 a_8327_3169.t3 a_8327_3169.t4 337.399
R9238 a_8327_3169.t4 a_8327_3169.t5 298.839
R9239 a_8327_3169.n0 a_8327_3169.t3 280.405
R9240 a_8327_3169.n1 a_8327_3169.t2 200
R9241 a_8327_3169.n1 a_8327_3169.n0 172.311
R9242 a_8327_3169.n2 a_8327_3169.n1 24
R9243 a_8327_3169.n1 a_8327_3169.t0 21.212
R9244 a_8422_3184.n0 a_8422_3184.t1 358.166
R9245 a_8422_3184.t5 a_8422_3184.t4 337.399
R9246 a_8422_3184.t4 a_8422_3184.t3 285.986
R9247 a_8422_3184.n0 a_8422_3184.t5 282.573
R9248 a_8422_3184.n1 a_8422_3184.t2 202.857
R9249 a_8422_3184.n1 a_8422_3184.n0 173.817
R9250 a_8422_3184.n1 a_8422_3184.t0 20.826
R9251 a_8422_3184.n2 a_8422_3184.n1 20.689
R9252 a_3152_2165.n0 a_3152_2165.t0 362.857
R9253 a_3152_2165.t3 a_3152_2165.t4 337.399
R9254 a_3152_2165.t4 a_3152_2165.t5 298.839
R9255 a_3152_2165.n0 a_3152_2165.t3 280.405
R9256 a_3152_2165.n1 a_3152_2165.t2 200
R9257 a_3152_2165.n1 a_3152_2165.n0 172.311
R9258 a_3152_2165.n2 a_3152_2165.n1 24
R9259 a_3152_2165.n1 a_3152_2165.t1 21.212
R9260 a_3247_2180.n0 a_3247_2180.t1 358.166
R9261 a_3247_2180.t4 a_3247_2180.t5 337.399
R9262 a_3247_2180.t5 a_3247_2180.t3 285.986
R9263 a_3247_2180.n0 a_3247_2180.t4 282.573
R9264 a_3247_2180.n1 a_3247_2180.t2 202.857
R9265 a_3247_2180.n1 a_3247_2180.n0 173.817
R9266 a_3247_2180.n1 a_3247_2180.t0 20.826
R9267 a_3247_2180.n2 a_3247_2180.n1 20.689
R9268 a_2035_n1371.n1 a_2035_n1371.t4 550.94
R9269 a_2035_n1371.n1 a_2035_n1371.t3 500.621
R9270 a_2035_n1371.t1 a_2035_n1371.n2 192.787
R9271 a_2035_n1371.n0 a_2035_n1371.t2 163.997
R9272 a_2035_n1371.n2 a_2035_n1371.n1 149.035
R9273 a_2035_n1371.n0 a_2035_n1371.t0 54.068
R9274 a_2035_n1371.n2 a_2035_n1371.n0 17.317
R9275 a_865_n812.t0 a_865_n812.t1 242.857
R9276 a_865_n953.t33 a_865_n953.n46 172.62
R9277 a_865_n953.n22 a_865_n953.t11 67.378
R9278 a_865_n953.n0 a_865_n953.t8 66.92
R9279 a_865_n953.n1 a_865_n953.t6 66.92
R9280 a_865_n953.n2 a_865_n953.t15 66.92
R9281 a_865_n953.n3 a_865_n953.t9 66.92
R9282 a_865_n953.n4 a_865_n953.t4 66.92
R9283 a_865_n953.n5 a_865_n953.t46 66.92
R9284 a_865_n953.n6 a_865_n953.t38 66.92
R9285 a_865_n953.n7 a_865_n953.t42 66.92
R9286 a_865_n953.n8 a_865_n953.t25 66.92
R9287 a_865_n953.n9 a_865_n953.t2 66.92
R9288 a_865_n953.n10 a_865_n953.t21 66.92
R9289 a_865_n953.n11 a_865_n953.t29 66.92
R9290 a_865_n953.n12 a_865_n953.t27 66.92
R9291 a_865_n953.n13 a_865_n953.t43 66.92
R9292 a_865_n953.n14 a_865_n953.t45 66.92
R9293 a_865_n953.n15 a_865_n953.t44 66.92
R9294 a_865_n953.n16 a_865_n953.t40 66.92
R9295 a_865_n953.n17 a_865_n953.t0 66.92
R9296 a_865_n953.n18 a_865_n953.t24 66.92
R9297 a_865_n953.n19 a_865_n953.t1 66.92
R9298 a_865_n953.n20 a_865_n953.t10 66.92
R9299 a_865_n953.n21 a_865_n953.t16 66.92
R9300 a_865_n953.n22 a_865_n953.t20 66.92
R9301 a_865_n953.n23 a_865_n953.t7 65.518
R9302 a_865_n953.n45 a_865_n953.t17 63.519
R9303 a_865_n953.n44 a_865_n953.t14 63.519
R9304 a_865_n953.n43 a_865_n953.t5 63.519
R9305 a_865_n953.n42 a_865_n953.t13 63.519
R9306 a_865_n953.n41 a_865_n953.t34 63.519
R9307 a_865_n953.n40 a_865_n953.t37 63.519
R9308 a_865_n953.n39 a_865_n953.t23 63.519
R9309 a_865_n953.n38 a_865_n953.t22 63.519
R9310 a_865_n953.n37 a_865_n953.t41 63.519
R9311 a_865_n953.n36 a_865_n953.t36 63.519
R9312 a_865_n953.n35 a_865_n953.t28 63.519
R9313 a_865_n953.n34 a_865_n953.t30 63.519
R9314 a_865_n953.n33 a_865_n953.t31 63.519
R9315 a_865_n953.n32 a_865_n953.t39 63.519
R9316 a_865_n953.n31 a_865_n953.t47 63.519
R9317 a_865_n953.n30 a_865_n953.t35 63.519
R9318 a_865_n953.n29 a_865_n953.t32 63.519
R9319 a_865_n953.n28 a_865_n953.t48 63.519
R9320 a_865_n953.n27 a_865_n953.t3 63.519
R9321 a_865_n953.n26 a_865_n953.t26 63.519
R9322 a_865_n953.n25 a_865_n953.t12 63.519
R9323 a_865_n953.n24 a_865_n953.t19 63.519
R9324 a_865_n953.n23 a_865_n953.t18 63.519
R9325 a_865_n953.n46 a_865_n953.n45 18.144
R9326 a_865_n953.n46 a_865_n953.n0 17.125
R9327 a_865_n953.n44 a_865_n953.n43 2.524
R9328 a_865_n953.n24 a_865_n953.n23 2.498
R9329 a_865_n953.n21 a_865_n953.n22 2.495
R9330 a_865_n953.n1 a_865_n953.n2 2.459
R9331 a_865_n953.n38 a_865_n953.n37 2.364
R9332 a_865_n953.n30 a_865_n953.n29 2.355
R9333 a_865_n953.n7 a_865_n953.n8 2.299
R9334 a_865_n953.n15 a_865_n953.n16 2.29
R9335 a_865_n953.n16 a_865_n953.n17 2.057
R9336 a_865_n953.n8 a_865_n953.n9 2.057
R9337 a_865_n953.n2 a_865_n953.n3 2.057
R9338 a_865_n953.n0 a_865_n953.n1 2.057
R9339 a_865_n953.n45 a_865_n953.n44 1.998
R9340 a_865_n953.n43 a_865_n953.n42 1.998
R9341 a_865_n953.n42 a_865_n953.n41 1.998
R9342 a_865_n953.n41 a_865_n953.n40 1.998
R9343 a_865_n953.n40 a_865_n953.n39 1.998
R9344 a_865_n953.n39 a_865_n953.n38 1.998
R9345 a_865_n953.n37 a_865_n953.n36 1.998
R9346 a_865_n953.n36 a_865_n953.n35 1.998
R9347 a_865_n953.n35 a_865_n953.n34 1.998
R9348 a_865_n953.n34 a_865_n953.n33 1.998
R9349 a_865_n953.n33 a_865_n953.n32 1.998
R9350 a_865_n953.n32 a_865_n953.n31 1.998
R9351 a_865_n953.n31 a_865_n953.n30 1.998
R9352 a_865_n953.n29 a_865_n953.n28 1.998
R9353 a_865_n953.n28 a_865_n953.n27 1.998
R9354 a_865_n953.n27 a_865_n953.n26 1.998
R9355 a_865_n953.n26 a_865_n953.n25 1.998
R9356 a_865_n953.n25 a_865_n953.n24 1.998
R9357 a_865_n953.n20 a_865_n953.n21 1.995
R9358 a_865_n953.n19 a_865_n953.n20 1.995
R9359 a_865_n953.n18 a_865_n953.n19 1.995
R9360 a_865_n953.n17 a_865_n953.n18 1.995
R9361 a_865_n953.n14 a_865_n953.n15 1.995
R9362 a_865_n953.n13 a_865_n953.n14 1.995
R9363 a_865_n953.n12 a_865_n953.n13 1.995
R9364 a_865_n953.n11 a_865_n953.n12 1.995
R9365 a_865_n953.n10 a_865_n953.n11 1.995
R9366 a_865_n953.n9 a_865_n953.n10 1.995
R9367 a_865_n953.n6 a_865_n953.n7 1.995
R9368 a_865_n953.n5 a_865_n953.n6 1.995
R9369 a_865_n953.n4 a_865_n953.n5 1.995
R9370 a_865_n953.n3 a_865_n953.n4 1.995
R9371 a_3740_4686.t0 a_3740_4686.t1 242.857
R9372 a_3740_n953.t34 a_3740_n953.n46 176.385
R9373 a_3740_n953.n22 a_3740_n953.t9 67.378
R9374 a_3740_n953.n0 a_3740_n953.t15 66.92
R9375 a_3740_n953.n1 a_3740_n953.t14 66.92
R9376 a_3740_n953.n2 a_3740_n953.t17 66.92
R9377 a_3740_n953.n3 a_3740_n953.t21 66.92
R9378 a_3740_n953.n4 a_3740_n953.t5 66.92
R9379 a_3740_n953.n5 a_3740_n953.t47 66.92
R9380 a_3740_n953.n6 a_3740_n953.t39 66.92
R9381 a_3740_n953.n7 a_3740_n953.t43 66.92
R9382 a_3740_n953.n8 a_3740_n953.t26 66.92
R9383 a_3740_n953.n9 a_3740_n953.t2 66.92
R9384 a_3740_n953.n10 a_3740_n953.t22 66.92
R9385 a_3740_n953.n11 a_3740_n953.t31 66.92
R9386 a_3740_n953.n12 a_3740_n953.t29 66.92
R9387 a_3740_n953.n13 a_3740_n953.t44 66.92
R9388 a_3740_n953.n14 a_3740_n953.t46 66.92
R9389 a_3740_n953.n15 a_3740_n953.t45 66.92
R9390 a_3740_n953.n16 a_3740_n953.t41 66.92
R9391 a_3740_n953.n17 a_3740_n953.t1 66.92
R9392 a_3740_n953.n18 a_3740_n953.t24 66.92
R9393 a_3740_n953.n19 a_3740_n953.t0 66.92
R9394 a_3740_n953.n20 a_3740_n953.t11 66.92
R9395 a_3740_n953.n21 a_3740_n953.t8 66.92
R9396 a_3740_n953.n22 a_3740_n953.t12 66.92
R9397 a_3740_n953.n23 a_3740_n953.t6 65.518
R9398 a_3740_n953.n45 a_3740_n953.t19 63.519
R9399 a_3740_n953.n44 a_3740_n953.t16 63.519
R9400 a_3740_n953.n43 a_3740_n953.t13 63.519
R9401 a_3740_n953.n42 a_3740_n953.t20 63.519
R9402 a_3740_n953.n41 a_3740_n953.t35 63.519
R9403 a_3740_n953.n40 a_3740_n953.t38 63.519
R9404 a_3740_n953.n39 a_3740_n953.t25 63.519
R9405 a_3740_n953.n38 a_3740_n953.t23 63.519
R9406 a_3740_n953.n37 a_3740_n953.t42 63.519
R9407 a_3740_n953.n36 a_3740_n953.t37 63.519
R9408 a_3740_n953.n35 a_3740_n953.t30 63.519
R9409 a_3740_n953.n34 a_3740_n953.t32 63.519
R9410 a_3740_n953.n33 a_3740_n953.t27 63.519
R9411 a_3740_n953.n32 a_3740_n953.t40 63.519
R9412 a_3740_n953.n31 a_3740_n953.t48 63.519
R9413 a_3740_n953.n30 a_3740_n953.t36 63.519
R9414 a_3740_n953.n29 a_3740_n953.t33 63.519
R9415 a_3740_n953.n28 a_3740_n953.t4 63.519
R9416 a_3740_n953.n27 a_3740_n953.t3 63.519
R9417 a_3740_n953.n26 a_3740_n953.t28 63.519
R9418 a_3740_n953.n25 a_3740_n953.t10 63.519
R9419 a_3740_n953.n24 a_3740_n953.t18 63.519
R9420 a_3740_n953.n23 a_3740_n953.t7 63.519
R9421 a_3740_n953.n46 a_3740_n953.n0 19.599
R9422 a_3740_n953.n46 a_3740_n953.n45 15.67
R9423 a_3740_n953.n44 a_3740_n953.n43 2.524
R9424 a_3740_n953.n24 a_3740_n953.n23 2.498
R9425 a_3740_n953.n21 a_3740_n953.n22 2.495
R9426 a_3740_n953.n1 a_3740_n953.n2 2.459
R9427 a_3740_n953.n38 a_3740_n953.n37 2.364
R9428 a_3740_n953.n30 a_3740_n953.n29 2.355
R9429 a_3740_n953.n7 a_3740_n953.n8 2.299
R9430 a_3740_n953.n15 a_3740_n953.n16 2.29
R9431 a_3740_n953.n16 a_3740_n953.n17 2.057
R9432 a_3740_n953.n8 a_3740_n953.n9 2.057
R9433 a_3740_n953.n2 a_3740_n953.n3 2.057
R9434 a_3740_n953.n0 a_3740_n953.n1 2.057
R9435 a_3740_n953.n45 a_3740_n953.n44 1.998
R9436 a_3740_n953.n43 a_3740_n953.n42 1.998
R9437 a_3740_n953.n42 a_3740_n953.n41 1.998
R9438 a_3740_n953.n41 a_3740_n953.n40 1.998
R9439 a_3740_n953.n40 a_3740_n953.n39 1.998
R9440 a_3740_n953.n39 a_3740_n953.n38 1.998
R9441 a_3740_n953.n37 a_3740_n953.n36 1.998
R9442 a_3740_n953.n36 a_3740_n953.n35 1.998
R9443 a_3740_n953.n35 a_3740_n953.n34 1.998
R9444 a_3740_n953.n34 a_3740_n953.n33 1.998
R9445 a_3740_n953.n33 a_3740_n953.n32 1.998
R9446 a_3740_n953.n32 a_3740_n953.n31 1.998
R9447 a_3740_n953.n31 a_3740_n953.n30 1.998
R9448 a_3740_n953.n29 a_3740_n953.n28 1.998
R9449 a_3740_n953.n28 a_3740_n953.n27 1.998
R9450 a_3740_n953.n27 a_3740_n953.n26 1.998
R9451 a_3740_n953.n26 a_3740_n953.n25 1.998
R9452 a_3740_n953.n25 a_3740_n953.n24 1.998
R9453 a_3740_n953.n20 a_3740_n953.n21 1.995
R9454 a_3740_n953.n19 a_3740_n953.n20 1.995
R9455 a_3740_n953.n18 a_3740_n953.n19 1.995
R9456 a_3740_n953.n17 a_3740_n953.n18 1.995
R9457 a_3740_n953.n14 a_3740_n953.n15 1.995
R9458 a_3740_n953.n13 a_3740_n953.n14 1.995
R9459 a_3740_n953.n12 a_3740_n953.n13 1.995
R9460 a_3740_n953.n11 a_3740_n953.n12 1.995
R9461 a_3740_n953.n10 a_3740_n953.n11 1.995
R9462 a_3740_n953.n9 a_3740_n953.n10 1.995
R9463 a_3740_n953.n6 a_3740_n953.n7 1.995
R9464 a_3740_n953.n5 a_3740_n953.n6 1.995
R9465 a_3740_n953.n4 a_3740_n953.n5 1.995
R9466 a_3740_n953.n3 a_3740_n953.n4 1.995
R9467 RWLB[1].n0 RWLB[1].t4 154.228
R9468 RWLB[1].n14 RWLB[1].t5 149.249
R9469 RWLB[1].n13 RWLB[1].t7 149.249
R9470 RWLB[1].n12 RWLB[1].t2 149.249
R9471 RWLB[1].n11 RWLB[1].t12 149.249
R9472 RWLB[1].n10 RWLB[1].t6 149.249
R9473 RWLB[1].n9 RWLB[1].t9 149.249
R9474 RWLB[1].n8 RWLB[1].t10 149.249
R9475 RWLB[1].n7 RWLB[1].t15 149.249
R9476 RWLB[1].n6 RWLB[1].t8 149.249
R9477 RWLB[1].n5 RWLB[1].t13 149.249
R9478 RWLB[1].n4 RWLB[1].t14 149.249
R9479 RWLB[1].n3 RWLB[1].t3 149.249
R9480 RWLB[1].n2 RWLB[1].t11 149.249
R9481 RWLB[1].n1 RWLB[1].t1 149.249
R9482 RWLB[1].n0 RWLB[1].t0 149.249
R9483 RWLB[1] RWLB[1].n14 47.816
R9484 RWLB[1].n1 RWLB[1].n0 4.979
R9485 RWLB[1].n2 RWLB[1].n1 4.979
R9486 RWLB[1].n3 RWLB[1].n2 4.979
R9487 RWLB[1].n4 RWLB[1].n3 4.979
R9488 RWLB[1].n5 RWLB[1].n4 4.979
R9489 RWLB[1].n6 RWLB[1].n5 4.979
R9490 RWLB[1].n7 RWLB[1].n6 4.979
R9491 RWLB[1].n8 RWLB[1].n7 4.979
R9492 RWLB[1].n9 RWLB[1].n8 4.979
R9493 RWLB[1].n10 RWLB[1].n9 4.979
R9494 RWLB[1].n11 RWLB[1].n10 4.979
R9495 RWLB[1].n12 RWLB[1].n11 4.979
R9496 RWLB[1].n13 RWLB[1].n12 4.979
R9497 RWLB[1].n14 RWLB[1].n13 4.979
R9498 a_8792_3425.t0 a_8792_3425.t1 242.857
R9499 a_4972_1698.n0 a_4972_1698.t0 358.166
R9500 a_4972_1698.t4 a_4972_1698.t3 337.399
R9501 a_4972_1698.t3 a_4972_1698.t5 285.986
R9502 a_4972_1698.n0 a_4972_1698.t4 282.573
R9503 a_4972_1698.n1 a_4972_1698.t2 202.857
R9504 a_4972_1698.n1 a_4972_1698.n0 173.817
R9505 a_4972_1698.n1 a_4972_1698.t1 20.826
R9506 a_4972_1698.n2 a_4972_1698.n1 20.689
R9507 a_4877_1683.n0 a_4877_1683.t1 362.857
R9508 a_4877_1683.t4 a_4877_1683.t3 337.399
R9509 a_4877_1683.t3 a_4877_1683.t5 298.839
R9510 a_4877_1683.n0 a_4877_1683.t4 280.405
R9511 a_4877_1683.n1 a_4877_1683.t2 200
R9512 a_4877_1683.n1 a_4877_1683.n0 172.311
R9513 a_4877_1683.n2 a_4877_1683.n1 24
R9514 a_4877_1683.n1 a_4877_1683.t0 21.212
R9515 a_8327_n45.n0 a_8327_n45.t0 362.857
R9516 a_8327_n45.t4 a_8327_n45.t3 337.399
R9517 a_8327_n45.t3 a_8327_n45.t5 298.839
R9518 a_8327_n45.n0 a_8327_n45.t4 280.405
R9519 a_8327_n45.n1 a_8327_n45.t2 200
R9520 a_8327_n45.n1 a_8327_n45.n0 172.311
R9521 a_8327_n45.n2 a_8327_n45.n1 24
R9522 a_8327_n45.n1 a_8327_n45.t1 21.212
R9523 a_8422_n30.n0 a_8422_n30.t1 358.166
R9524 a_8422_n30.t5 a_8422_n30.t3 337.399
R9525 a_8422_n30.t3 a_8422_n30.t4 285.986
R9526 a_8422_n30.n0 a_8422_n30.t5 282.573
R9527 a_8422_n30.n1 a_8422_n30.t2 202.857
R9528 a_8422_n30.n1 a_8422_n30.n0 173.817
R9529 a_8422_n30.n1 a_8422_n30.t0 20.826
R9530 a_8422_n30.n2 a_8422_n30.n1 20.689
R9531 ADC10_OUT[2].n0 ADC10_OUT[2].t4 1354.27
R9532 ADC10_OUT[2].n0 ADC10_OUT[2].t3 821.954
R9533 ADC10_OUT[2].n3 ADC10_OUT[2].t2 338.103
R9534 ADC10_OUT[2].n2 ADC10_OUT[2].t0 266.575
R9535 ADC10_OUT[2].n1 ADC10_OUT[2].n0 149.035
R9536 ADC10_OUT[2].n1 ADC10_OUT[2].t1 46.723
R9537 ADC10_OUT[2].n3 ADC10_OUT[2].n2 45.929
R9538 ADC10_OUT[2] ADC10_OUT[2].n3 38.172
R9539 ADC10_OUT[2].n2 ADC10_OUT[2].n1 17.317
R9540 a_8221_n7216.n0 a_8221_n7216.t3 1464.36
R9541 a_8221_n7216.n0 a_8221_n7216.t4 713.588
R9542 a_8221_n7216.n1 a_8221_n7216.t0 374.998
R9543 a_8221_n7216.n1 a_8221_n7216.t1 273.351
R9544 a_8221_n7216.n2 a_8221_n7216.n0 143.764
R9545 a_8221_n7216.t2 a_8221_n7216.n2 78.209
R9546 a_8221_n7216.n2 a_8221_n7216.n1 4.517
R9547 a_4397_n812.n0 a_4397_n812.t1 358.166
R9548 a_4397_n812.t4 a_4397_n812.t5 337.399
R9549 a_4397_n812.t5 a_4397_n812.t3 285.986
R9550 a_4397_n812.n0 a_4397_n812.t4 282.573
R9551 a_4397_n812.n1 a_4397_n812.t0 202.857
R9552 a_4397_n812.n1 a_4397_n812.n0 173.817
R9553 a_4397_n812.n1 a_4397_n812.t2 20.826
R9554 a_4397_n812.n2 a_4397_n812.n1 20.689
R9555 a_4767_n812.t0 a_4767_n812.t1 242.857
R9556 WWL[1].n0 WWL[1].t6 262.032
R9557 WWL[1].n29 WWL[1].t9 260.715
R9558 WWL[1].n27 WWL[1].t12 260.715
R9559 WWL[1].n25 WWL[1].t26 260.715
R9560 WWL[1].n23 WWL[1].t20 260.715
R9561 WWL[1].n21 WWL[1].t0 260.715
R9562 WWL[1].n19 WWL[1].t17 260.715
R9563 WWL[1].n17 WWL[1].t8 260.715
R9564 WWL[1].n15 WWL[1].t23 260.715
R9565 WWL[1].n13 WWL[1].t13 260.715
R9566 WWL[1].n11 WWL[1].t21 260.715
R9567 WWL[1].n9 WWL[1].t10 260.715
R9568 WWL[1].n7 WWL[1].t24 260.715
R9569 WWL[1].n5 WWL[1].t18 260.715
R9570 WWL[1].n3 WWL[1].t1 260.715
R9571 WWL[1].n1 WWL[1].t14 260.715
R9572 WWL[1].n30 WWL[1].t25 259.254
R9573 WWL[1].n28 WWL[1].t31 259.254
R9574 WWL[1].n26 WWL[1].t11 259.254
R9575 WWL[1].n24 WWL[1].t27 259.254
R9576 WWL[1].n22 WWL[1].t19 259.254
R9577 WWL[1].n20 WWL[1].t2 259.254
R9578 WWL[1].n18 WWL[1].t15 259.254
R9579 WWL[1].n16 WWL[1].t29 259.254
R9580 WWL[1].n14 WWL[1].t22 259.254
R9581 WWL[1].n12 WWL[1].t5 259.254
R9582 WWL[1].n10 WWL[1].t28 259.254
R9583 WWL[1].n8 WWL[1].t3 259.254
R9584 WWL[1].n6 WWL[1].t4 259.254
R9585 WWL[1].n4 WWL[1].t7 259.254
R9586 WWL[1].n2 WWL[1].t30 259.254
R9587 WWL[1].n0 WWL[1].t16 259.254
R9588 WWL[1] WWL[1].n30 44.647
R9589 WWL[1].n1 WWL[1].n0 3.576
R9590 WWL[1].n3 WWL[1].n2 3.576
R9591 WWL[1].n5 WWL[1].n4 3.576
R9592 WWL[1].n7 WWL[1].n6 3.576
R9593 WWL[1].n9 WWL[1].n8 3.576
R9594 WWL[1].n11 WWL[1].n10 3.576
R9595 WWL[1].n13 WWL[1].n12 3.576
R9596 WWL[1].n15 WWL[1].n14 3.576
R9597 WWL[1].n17 WWL[1].n16 3.576
R9598 WWL[1].n19 WWL[1].n18 3.576
R9599 WWL[1].n21 WWL[1].n20 3.576
R9600 WWL[1].n23 WWL[1].n22 3.576
R9601 WWL[1].n25 WWL[1].n24 3.576
R9602 WWL[1].n27 WWL[1].n26 3.576
R9603 WWL[1].n29 WWL[1].n28 3.576
R9604 WWL[1].n2 WWL[1].n1 1.317
R9605 WWL[1].n4 WWL[1].n3 1.317
R9606 WWL[1].n6 WWL[1].n5 1.317
R9607 WWL[1].n8 WWL[1].n7 1.317
R9608 WWL[1].n10 WWL[1].n9 1.317
R9609 WWL[1].n12 WWL[1].n11 1.317
R9610 WWL[1].n14 WWL[1].n13 1.317
R9611 WWL[1].n16 WWL[1].n15 1.317
R9612 WWL[1].n18 WWL[1].n17 1.317
R9613 WWL[1].n20 WWL[1].n19 1.317
R9614 WWL[1].n22 WWL[1].n21 1.317
R9615 WWL[1].n24 WWL[1].n23 1.317
R9616 WWL[1].n26 WWL[1].n25 1.317
R9617 WWL[1].n28 WWL[1].n27 1.317
R9618 WWL[1].n30 WWL[1].n29 1.317
R9619 a_2845_4887.n25 a_2845_4887.t27 561.971
R9620 a_2845_4887.n0 a_2845_4887.t19 449.944
R9621 a_2845_4887.t26 a_2845_4887.n25 108.636
R9622 a_2845_4887.n0 a_2845_4887.t20 74.821
R9623 a_2845_4887.n24 a_2845_4887.t23 63.519
R9624 a_2845_4887.n23 a_2845_4887.t6 63.519
R9625 a_2845_4887.n22 a_2845_4887.t5 63.519
R9626 a_2845_4887.n21 a_2845_4887.t16 63.519
R9627 a_2845_4887.n20 a_2845_4887.t9 63.519
R9628 a_2845_4887.n19 a_2845_4887.t17 63.519
R9629 a_2845_4887.n18 a_2845_4887.t22 63.519
R9630 a_2845_4887.n17 a_2845_4887.t14 63.519
R9631 a_2845_4887.n16 a_2845_4887.t21 63.519
R9632 a_2845_4887.n15 a_2845_4887.t2 63.519
R9633 a_2845_4887.n14 a_2845_4887.t13 63.519
R9634 a_2845_4887.n13 a_2845_4887.t10 63.519
R9635 a_2845_4887.n12 a_2845_4887.t1 63.519
R9636 a_2845_4887.n11 a_2845_4887.t12 63.519
R9637 a_2845_4887.n10 a_2845_4887.t4 63.519
R9638 a_2845_4887.n9 a_2845_4887.t8 63.519
R9639 a_2845_4887.n8 a_2845_4887.t7 63.519
R9640 a_2845_4887.n7 a_2845_4887.t24 63.519
R9641 a_2845_4887.n6 a_2845_4887.t3 63.519
R9642 a_2845_4887.n5 a_2845_4887.t25 63.519
R9643 a_2845_4887.n4 a_2845_4887.t0 63.519
R9644 a_2845_4887.n3 a_2845_4887.t11 63.519
R9645 a_2845_4887.n2 a_2845_4887.t15 63.519
R9646 a_2845_4887.n1 a_2845_4887.t18 63.519
R9647 a_2845_4887.n1 a_2845_4887.n0 8.619
R9648 a_2845_4887.n25 a_2845_4887.n24 2.946
R9649 a_2845_4887.n23 a_2845_4887.n22 2.524
R9650 a_2845_4887.n3 a_2845_4887.n2 2.498
R9651 a_2845_4887.n17 a_2845_4887.n16 2.364
R9652 a_2845_4887.n9 a_2845_4887.n8 2.355
R9653 a_2845_4887.n24 a_2845_4887.n23 1.998
R9654 a_2845_4887.n22 a_2845_4887.n21 1.998
R9655 a_2845_4887.n21 a_2845_4887.n20 1.998
R9656 a_2845_4887.n20 a_2845_4887.n19 1.998
R9657 a_2845_4887.n19 a_2845_4887.n18 1.998
R9658 a_2845_4887.n18 a_2845_4887.n17 1.998
R9659 a_2845_4887.n16 a_2845_4887.n15 1.998
R9660 a_2845_4887.n15 a_2845_4887.n14 1.998
R9661 a_2845_4887.n14 a_2845_4887.n13 1.998
R9662 a_2845_4887.n13 a_2845_4887.n12 1.998
R9663 a_2845_4887.n12 a_2845_4887.n11 1.998
R9664 a_2845_4887.n11 a_2845_4887.n10 1.998
R9665 a_2845_4887.n10 a_2845_4887.n9 1.998
R9666 a_2845_4887.n8 a_2845_4887.n7 1.998
R9667 a_2845_4887.n7 a_2845_4887.n6 1.998
R9668 a_2845_4887.n6 a_2845_4887.n5 1.998
R9669 a_2845_4887.n5 a_2845_4887.n4 1.998
R9670 a_2845_4887.n4 a_2845_4887.n3 1.998
R9671 a_2845_4887.n2 a_2845_4887.n1 1.998
R9672 a_2577_3410.n0 a_2577_3410.t2 362.857
R9673 a_2577_3410.t3 a_2577_3410.t4 337.399
R9674 a_2577_3410.t4 a_2577_3410.t5 298.839
R9675 a_2577_3410.n0 a_2577_3410.t3 280.405
R9676 a_2577_3410.n1 a_2577_3410.t0 200
R9677 a_2577_3410.n1 a_2577_3410.n0 172.311
R9678 a_2577_3410.n2 a_2577_3410.n1 24
R9679 a_2577_3410.n1 a_2577_3410.t1 21.212
R9680 a_3727_678.n0 a_3727_678.t0 362.857
R9681 a_3727_678.t3 a_3727_678.t5 337.399
R9682 a_3727_678.t5 a_3727_678.t4 298.839
R9683 a_3727_678.n0 a_3727_678.t3 280.405
R9684 a_3727_678.n1 a_3727_678.t2 200
R9685 a_3727_678.n1 a_3727_678.n0 172.311
R9686 a_3727_678.n2 a_3727_678.n1 24
R9687 a_3727_678.n1 a_3727_678.t1 21.212
R9688 a_3822_693.n0 a_3822_693.t1 358.166
R9689 a_3822_693.t3 a_3822_693.t5 337.399
R9690 a_3822_693.t5 a_3822_693.t4 285.986
R9691 a_3822_693.n0 a_3822_693.t3 282.573
R9692 a_3822_693.n1 a_3822_693.t2 202.857
R9693 a_3822_693.n1 a_3822_693.n0 173.817
R9694 a_3822_693.n1 a_3822_693.t0 20.826
R9695 a_3822_693.n2 a_3822_693.n1 20.689
R9696 SAEN.n63 SAEN.t21 187.425
R9697 SAEN.n0 SAEN.t55 187.425
R9698 SAEN.n77 SAEN.t6 186.057
R9699 SAEN.n75 SAEN.t42 186.057
R9700 SAEN.n73 SAEN.t92 186.057
R9701 SAEN.n71 SAEN.t81 186.057
R9702 SAEN.n69 SAEN.t34 186.057
R9703 SAEN.n67 SAEN.t74 186.057
R9704 SAEN.n65 SAEN.t111 186.057
R9705 SAEN.n63 SAEN.t79 186.057
R9706 SAEN.n30 SAEN.t10 186.057
R9707 SAEN.n28 SAEN.t50 186.057
R9708 SAEN.n26 SAEN.t95 186.057
R9709 SAEN.n24 SAEN.t84 186.057
R9710 SAEN.n22 SAEN.t38 186.057
R9711 SAEN.n20 SAEN.t78 186.057
R9712 SAEN.n18 SAEN.t1 186.057
R9713 SAEN.n16 SAEN.t82 186.057
R9714 SAEN.n14 SAEN.t31 186.057
R9715 SAEN.n12 SAEN.t4 186.057
R9716 SAEN.n10 SAEN.t33 186.057
R9717 SAEN.n8 SAEN.t48 186.057
R9718 SAEN.n6 SAEN.t36 186.057
R9719 SAEN.n4 SAEN.t30 186.057
R9720 SAEN.n2 SAEN.t23 186.057
R9721 SAEN.n0 SAEN.t2 186.057
R9722 SAEN.n79 SAEN.t32 184.212
R9723 SAEN.n31 SAEN.t83 184.212
R9724 SAEN.n109 SAEN.t0 182.844
R9725 SAEN.n107 SAEN.t29 182.844
R9726 SAEN.n105 SAEN.t73 182.844
R9727 SAEN.n103 SAEN.t61 182.844
R9728 SAEN.n101 SAEN.t22 182.844
R9729 SAEN.n99 SAEN.t52 182.844
R9730 SAEN.n97 SAEN.t100 182.844
R9731 SAEN.n95 SAEN.t56 182.844
R9732 SAEN.n93 SAEN.t15 182.844
R9733 SAEN.n91 SAEN.t106 182.844
R9734 SAEN.n89 SAEN.t16 182.844
R9735 SAEN.n87 SAEN.t26 182.844
R9736 SAEN.n85 SAEN.t19 182.844
R9737 SAEN.n83 SAEN.t13 182.844
R9738 SAEN.n81 SAEN.t7 182.844
R9739 SAEN.n79 SAEN.t105 182.844
R9740 SAEN.n61 SAEN.t27 182.844
R9741 SAEN.n59 SAEN.t77 182.844
R9742 SAEN.n57 SAEN.t109 182.844
R9743 SAEN.n55 SAEN.t103 182.844
R9744 SAEN.n53 SAEN.t67 182.844
R9745 SAEN.n51 SAEN.t97 182.844
R9746 SAEN.n49 SAEN.t12 182.844
R9747 SAEN.n47 SAEN.t101 182.844
R9748 SAEN.n45 SAEN.t58 182.844
R9749 SAEN.n43 SAEN.t18 182.844
R9750 SAEN.n41 SAEN.t60 182.844
R9751 SAEN.n39 SAEN.t72 182.844
R9752 SAEN.n37 SAEN.t66 182.844
R9753 SAEN.n35 SAEN.t51 182.844
R9754 SAEN.n33 SAEN.t44 182.844
R9755 SAEN.n31 SAEN.t14 182.844
R9756 SAEN.n76 SAEN.t54 182.843
R9757 SAEN.n74 SAEN.t99 182.843
R9758 SAEN.n72 SAEN.t41 182.843
R9759 SAEN.n70 SAEN.t75 182.843
R9760 SAEN.n68 SAEN.t57 182.843
R9761 SAEN.n66 SAEN.t17 182.843
R9762 SAEN.n64 SAEN.t65 182.843
R9763 SAEN.n29 SAEN.t59 182.843
R9764 SAEN.n27 SAEN.t102 182.843
R9765 SAEN.n25 SAEN.t49 182.843
R9766 SAEN.n23 SAEN.t80 182.843
R9767 SAEN.n21 SAEN.t64 182.843
R9768 SAEN.n19 SAEN.t20 182.843
R9769 SAEN.n17 SAEN.t69 182.843
R9770 SAEN.n15 SAEN.t24 182.843
R9771 SAEN.n13 SAEN.t70 182.843
R9772 SAEN.n11 SAEN.t25 182.843
R9773 SAEN.n9 SAEN.t110 182.843
R9774 SAEN.n7 SAEN.t85 182.843
R9775 SAEN.n5 SAEN.t89 182.843
R9776 SAEN.n3 SAEN.t63 182.843
R9777 SAEN.n1 SAEN.t91 182.843
R9778 SAEN.n108 SAEN.t35 179.63
R9779 SAEN.n106 SAEN.t87 179.63
R9780 SAEN.n104 SAEN.t28 179.63
R9781 SAEN.n102 SAEN.t53 179.63
R9782 SAEN.n100 SAEN.t39 179.63
R9783 SAEN.n98 SAEN.t5 179.63
R9784 SAEN.n96 SAEN.t43 179.63
R9785 SAEN.n94 SAEN.t8 179.63
R9786 SAEN.n92 SAEN.t45 179.63
R9787 SAEN.n90 SAEN.t9 179.63
R9788 SAEN.n88 SAEN.t96 179.63
R9789 SAEN.n86 SAEN.t62 179.63
R9790 SAEN.n84 SAEN.t68 179.63
R9791 SAEN.n82 SAEN.t37 179.63
R9792 SAEN.n80 SAEN.t71 179.63
R9793 SAEN.n60 SAEN.t86 179.63
R9794 SAEN.n58 SAEN.t3 179.63
R9795 SAEN.n56 SAEN.t76 179.63
R9796 SAEN.n54 SAEN.t98 179.63
R9797 SAEN.n52 SAEN.t90 179.63
R9798 SAEN.n50 SAEN.t40 179.63
R9799 SAEN.n48 SAEN.t93 179.63
R9800 SAEN.n46 SAEN.t46 179.63
R9801 SAEN.n44 SAEN.t94 179.63
R9802 SAEN.n42 SAEN.t47 179.63
R9803 SAEN.n40 SAEN.t11 179.63
R9804 SAEN.n38 SAEN.t104 179.63
R9805 SAEN.n36 SAEN.t107 179.63
R9806 SAEN.n34 SAEN.t88 179.63
R9807 SAEN.n32 SAEN.t108 179.63
R9808 SAEN.n62 SAEN.n30 21.895
R9809 SAEN.n110 SAEN.n78 14.534
R9810 SAEN.n78 SAEN.n62 9.543
R9811 SAEN SAEN.n110 8.526
R9812 SAEN.n110 SAEN.n109 7.347
R9813 SAEN.n78 SAEN.n77 7.347
R9814 SAEN.n62 SAEN.n61 7.347
R9815 SAEN.n82 SAEN.n81 5.78
R9816 SAEN.n84 SAEN.n83 5.78
R9817 SAEN.n34 SAEN.n33 5.78
R9818 SAEN.n36 SAEN.n35 5.78
R9819 SAEN.n3 SAEN.n2 5.78
R9820 SAEN.n5 SAEN.n4 5.78
R9821 SAEN.n86 SAEN.n85 5.753
R9822 SAEN.n88 SAEN.n87 5.753
R9823 SAEN.n38 SAEN.n37 5.753
R9824 SAEN.n40 SAEN.n39 5.753
R9825 SAEN.n7 SAEN.n6 5.753
R9826 SAEN.n9 SAEN.n8 5.753
R9827 SAEN.n90 SAEN.n89 5.735
R9828 SAEN.n92 SAEN.n91 5.735
R9829 SAEN.n94 SAEN.n93 5.735
R9830 SAEN.n96 SAEN.n95 5.735
R9831 SAEN.n98 SAEN.n97 5.735
R9832 SAEN.n100 SAEN.n99 5.735
R9833 SAEN.n106 SAEN.n105 5.735
R9834 SAEN.n64 SAEN.n63 5.735
R9835 SAEN.n66 SAEN.n65 5.735
R9836 SAEN.n68 SAEN.n67 5.735
R9837 SAEN.n74 SAEN.n73 5.735
R9838 SAEN.n42 SAEN.n41 5.735
R9839 SAEN.n44 SAEN.n43 5.735
R9840 SAEN.n46 SAEN.n45 5.735
R9841 SAEN.n48 SAEN.n47 5.735
R9842 SAEN.n50 SAEN.n49 5.735
R9843 SAEN.n52 SAEN.n51 5.735
R9844 SAEN.n58 SAEN.n57 5.735
R9845 SAEN.n11 SAEN.n10 5.735
R9846 SAEN.n13 SAEN.n12 5.735
R9847 SAEN.n15 SAEN.n14 5.735
R9848 SAEN.n17 SAEN.n16 5.735
R9849 SAEN.n19 SAEN.n18 5.735
R9850 SAEN.n21 SAEN.n20 5.735
R9851 SAEN.n27 SAEN.n26 5.735
R9852 SAEN.n102 SAEN.n101 5.726
R9853 SAEN.n104 SAEN.n103 5.726
R9854 SAEN.n70 SAEN.n69 5.726
R9855 SAEN.n72 SAEN.n71 5.726
R9856 SAEN.n54 SAEN.n53 5.726
R9857 SAEN.n56 SAEN.n55 5.726
R9858 SAEN.n23 SAEN.n22 5.726
R9859 SAEN.n25 SAEN.n24 5.726
R9860 SAEN.n108 SAEN.n107 5.449
R9861 SAEN.n76 SAEN.n75 5.449
R9862 SAEN.n60 SAEN.n59 5.449
R9863 SAEN.n29 SAEN.n28 5.449
R9864 SAEN.n81 SAEN.n80 4.582
R9865 SAEN.n83 SAEN.n82 4.582
R9866 SAEN.n85 SAEN.n84 4.582
R9867 SAEN.n87 SAEN.n86 4.582
R9868 SAEN.n89 SAEN.n88 4.582
R9869 SAEN.n91 SAEN.n90 4.582
R9870 SAEN.n93 SAEN.n92 4.582
R9871 SAEN.n95 SAEN.n94 4.582
R9872 SAEN.n97 SAEN.n96 4.582
R9873 SAEN.n99 SAEN.n98 4.582
R9874 SAEN.n101 SAEN.n100 4.582
R9875 SAEN.n103 SAEN.n102 4.582
R9876 SAEN.n105 SAEN.n104 4.582
R9877 SAEN.n107 SAEN.n106 4.582
R9878 SAEN.n109 SAEN.n108 4.582
R9879 SAEN.n65 SAEN.n64 4.582
R9880 SAEN.n67 SAEN.n66 4.582
R9881 SAEN.n69 SAEN.n68 4.582
R9882 SAEN.n71 SAEN.n70 4.582
R9883 SAEN.n73 SAEN.n72 4.582
R9884 SAEN.n75 SAEN.n74 4.582
R9885 SAEN.n77 SAEN.n76 4.582
R9886 SAEN.n33 SAEN.n32 4.582
R9887 SAEN.n35 SAEN.n34 4.582
R9888 SAEN.n37 SAEN.n36 4.582
R9889 SAEN.n39 SAEN.n38 4.582
R9890 SAEN.n41 SAEN.n40 4.582
R9891 SAEN.n43 SAEN.n42 4.582
R9892 SAEN.n45 SAEN.n44 4.582
R9893 SAEN.n47 SAEN.n46 4.582
R9894 SAEN.n49 SAEN.n48 4.582
R9895 SAEN.n51 SAEN.n50 4.582
R9896 SAEN.n53 SAEN.n52 4.582
R9897 SAEN.n55 SAEN.n54 4.582
R9898 SAEN.n57 SAEN.n56 4.582
R9899 SAEN.n59 SAEN.n58 4.582
R9900 SAEN.n61 SAEN.n60 4.582
R9901 SAEN.n2 SAEN.n1 4.582
R9902 SAEN.n4 SAEN.n3 4.582
R9903 SAEN.n6 SAEN.n5 4.582
R9904 SAEN.n8 SAEN.n7 4.582
R9905 SAEN.n10 SAEN.n9 4.582
R9906 SAEN.n12 SAEN.n11 4.582
R9907 SAEN.n14 SAEN.n13 4.582
R9908 SAEN.n16 SAEN.n15 4.582
R9909 SAEN.n18 SAEN.n17 4.582
R9910 SAEN.n20 SAEN.n19 4.582
R9911 SAEN.n22 SAEN.n21 4.582
R9912 SAEN.n24 SAEN.n23 4.582
R9913 SAEN.n26 SAEN.n25 4.582
R9914 SAEN.n28 SAEN.n27 4.582
R9915 SAEN.n30 SAEN.n29 4.582
R9916 SAEN.n80 SAEN.n79 3.226
R9917 SAEN.n32 SAEN.n31 3.226
R9918 SAEN.n1 SAEN.n0 3.226
R9919 a_n3792_n8026.n0 a_n3792_n8026.t1 65.063
R9920 a_n3792_n8026.n0 a_n3792_n8026.t2 42.011
R9921 a_n3792_n8026.t0 a_n3792_n8026.n0 2.113
R9922 PRE_CLSA.n95 PRE_CLSA.t119 737.3
R9923 PRE_CLSA.n0 PRE_CLSA.t100 735.84
R9924 PRE_CLSA.n125 PRE_CLSA.t78 733.783
R9925 PRE_CLSA.n124 PRE_CLSA.t124 733.783
R9926 PRE_CLSA.n123 PRE_CLSA.t76 733.783
R9927 PRE_CLSA.n122 PRE_CLSA.t123 733.783
R9928 PRE_CLSA.n121 PRE_CLSA.t20 733.783
R9929 PRE_CLSA.n120 PRE_CLSA.t40 733.783
R9930 PRE_CLSA.n119 PRE_CLSA.t52 733.783
R9931 PRE_CLSA.n118 PRE_CLSA.t0 733.783
R9932 PRE_CLSA.n117 PRE_CLSA.t35 733.783
R9933 PRE_CLSA.n116 PRE_CLSA.t114 733.783
R9934 PRE_CLSA.n115 PRE_CLSA.t99 733.783
R9935 PRE_CLSA.n114 PRE_CLSA.t44 733.783
R9936 PRE_CLSA.n113 PRE_CLSA.t57 733.783
R9937 PRE_CLSA.n112 PRE_CLSA.t2 733.783
R9938 PRE_CLSA.n111 PRE_CLSA.t18 733.783
R9939 PRE_CLSA.n110 PRE_CLSA.t94 733.783
R9940 PRE_CLSA.n109 PRE_CLSA.t75 733.783
R9941 PRE_CLSA.n108 PRE_CLSA.t37 733.783
R9942 PRE_CLSA.n107 PRE_CLSA.t113 733.783
R9943 PRE_CLSA.n106 PRE_CLSA.t84 733.783
R9944 PRE_CLSA.n105 PRE_CLSA.t61 733.783
R9945 PRE_CLSA.n104 PRE_CLSA.t8 733.783
R9946 PRE_CLSA.n103 PRE_CLSA.t74 733.783
R9947 PRE_CLSA.n102 PRE_CLSA.t22 733.783
R9948 PRE_CLSA.n101 PRE_CLSA.t80 733.783
R9949 PRE_CLSA.n100 PRE_CLSA.t55 733.783
R9950 PRE_CLSA.n99 PRE_CLSA.t67 733.783
R9951 PRE_CLSA.n98 PRE_CLSA.t33 733.783
R9952 PRE_CLSA.n97 PRE_CLSA.t92 733.783
R9953 PRE_CLSA.n96 PRE_CLSA.t24 733.783
R9954 PRE_CLSA.n95 PRE_CLSA.t63 733.783
R9955 PRE_CLSA.n30 PRE_CLSA.t49 732.323
R9956 PRE_CLSA.n29 PRE_CLSA.t105 732.323
R9957 PRE_CLSA.n28 PRE_CLSA.t48 732.323
R9958 PRE_CLSA.n27 PRE_CLSA.t102 732.323
R9959 PRE_CLSA.n26 PRE_CLSA.t118 732.323
R9960 PRE_CLSA.n25 PRE_CLSA.t19 732.323
R9961 PRE_CLSA.n24 PRE_CLSA.t28 732.323
R9962 PRE_CLSA.n23 PRE_CLSA.t107 732.323
R9963 PRE_CLSA.n22 PRE_CLSA.t13 732.323
R9964 PRE_CLSA.n21 PRE_CLSA.t96 732.323
R9965 PRE_CLSA.n20 PRE_CLSA.t79 732.323
R9966 PRE_CLSA.n19 PRE_CLSA.t23 732.323
R9967 PRE_CLSA.n18 PRE_CLSA.t34 732.323
R9968 PRE_CLSA.n17 PRE_CLSA.t110 732.323
R9969 PRE_CLSA.n16 PRE_CLSA.t117 732.323
R9970 PRE_CLSA.n15 PRE_CLSA.t71 732.323
R9971 PRE_CLSA.n14 PRE_CLSA.t47 732.323
R9972 PRE_CLSA.n13 PRE_CLSA.t15 732.323
R9973 PRE_CLSA.n12 PRE_CLSA.t95 732.323
R9974 PRE_CLSA.n11 PRE_CLSA.t58 732.323
R9975 PRE_CLSA.n10 PRE_CLSA.t38 732.323
R9976 PRE_CLSA.n9 PRE_CLSA.t111 732.323
R9977 PRE_CLSA.n8 PRE_CLSA.t46 732.323
R9978 PRE_CLSA.n7 PRE_CLSA.t120 732.323
R9979 PRE_CLSA.n6 PRE_CLSA.t53 732.323
R9980 PRE_CLSA.n5 PRE_CLSA.t31 732.323
R9981 PRE_CLSA.n4 PRE_CLSA.t42 732.323
R9982 PRE_CLSA.n3 PRE_CLSA.t11 732.323
R9983 PRE_CLSA.n2 PRE_CLSA.t70 732.323
R9984 PRE_CLSA.n1 PRE_CLSA.t127 732.323
R9985 PRE_CLSA.n0 PRE_CLSA.t39 732.323
R9986 PRE_CLSA.n92 PRE_CLSA.t89 720.369
R9987 PRE_CLSA.n90 PRE_CLSA.t10 720.369
R9988 PRE_CLSA.n88 PRE_CLSA.t88 720.369
R9989 PRE_CLSA.n86 PRE_CLSA.t7 720.369
R9990 PRE_CLSA.n84 PRE_CLSA.t29 720.369
R9991 PRE_CLSA.n82 PRE_CLSA.t51 720.369
R9992 PRE_CLSA.n80 PRE_CLSA.t64 720.369
R9993 PRE_CLSA.n78 PRE_CLSA.t14 720.369
R9994 PRE_CLSA.n76 PRE_CLSA.t43 720.369
R9995 PRE_CLSA.n74 PRE_CLSA.t126 720.369
R9996 PRE_CLSA.n72 PRE_CLSA.t109 720.369
R9997 PRE_CLSA.n70 PRE_CLSA.t56 720.369
R9998 PRE_CLSA.n68 PRE_CLSA.t69 720.369
R9999 PRE_CLSA.n66 PRE_CLSA.t16 720.369
R10000 PRE_CLSA.n64 PRE_CLSA.t27 720.369
R10001 PRE_CLSA.n62 PRE_CLSA.t104 720.369
R10002 PRE_CLSA.n60 PRE_CLSA.t87 720.369
R10003 PRE_CLSA.n58 PRE_CLSA.t45 720.369
R10004 PRE_CLSA.n56 PRE_CLSA.t125 720.369
R10005 PRE_CLSA.n54 PRE_CLSA.t93 720.369
R10006 PRE_CLSA.n52 PRE_CLSA.t73 720.369
R10007 PRE_CLSA.n50 PRE_CLSA.t21 720.369
R10008 PRE_CLSA.n48 PRE_CLSA.t86 720.369
R10009 PRE_CLSA.n46 PRE_CLSA.t30 720.369
R10010 PRE_CLSA.n44 PRE_CLSA.t90 720.369
R10011 PRE_CLSA.n42 PRE_CLSA.t66 720.369
R10012 PRE_CLSA.n40 PRE_CLSA.t81 720.369
R10013 PRE_CLSA.n38 PRE_CLSA.t41 720.369
R10014 PRE_CLSA.n36 PRE_CLSA.t103 720.369
R10015 PRE_CLSA.n34 PRE_CLSA.t36 720.369
R10016 PRE_CLSA.n32 PRE_CLSA.t77 720.369
R10017 PRE_CLSA.n31 PRE_CLSA.t3 720.369
R10018 PRE_CLSA.n92 PRE_CLSA.t9 718.909
R10019 PRE_CLSA.n90 PRE_CLSA.t62 718.909
R10020 PRE_CLSA.n88 PRE_CLSA.t6 718.909
R10021 PRE_CLSA.n86 PRE_CLSA.t60 718.909
R10022 PRE_CLSA.n84 PRE_CLSA.t83 718.909
R10023 PRE_CLSA.n82 PRE_CLSA.t106 718.909
R10024 PRE_CLSA.n80 PRE_CLSA.t112 718.909
R10025 PRE_CLSA.n78 PRE_CLSA.t65 718.909
R10026 PRE_CLSA.n76 PRE_CLSA.t98 718.909
R10027 PRE_CLSA.n74 PRE_CLSA.t54 718.909
R10028 PRE_CLSA.n72 PRE_CLSA.t32 718.909
R10029 PRE_CLSA.n70 PRE_CLSA.t108 718.909
R10030 PRE_CLSA.n68 PRE_CLSA.t116 718.909
R10031 PRE_CLSA.n66 PRE_CLSA.t68 718.909
R10032 PRE_CLSA.n64 PRE_CLSA.t82 718.909
R10033 PRE_CLSA.n62 PRE_CLSA.t26 718.909
R10034 PRE_CLSA.n60 PRE_CLSA.t5 718.909
R10035 PRE_CLSA.n58 PRE_CLSA.t101 718.909
R10036 PRE_CLSA.n56 PRE_CLSA.t50 718.909
R10037 PRE_CLSA.n54 PRE_CLSA.t17 718.909
R10038 PRE_CLSA.n52 PRE_CLSA.t121 718.909
R10039 PRE_CLSA.n50 PRE_CLSA.t72 718.909
R10040 PRE_CLSA.n48 PRE_CLSA.t4 718.909
R10041 PRE_CLSA.n46 PRE_CLSA.t85 718.909
R10042 PRE_CLSA.n44 PRE_CLSA.t12 718.909
R10043 PRE_CLSA.n42 PRE_CLSA.t115 718.909
R10044 PRE_CLSA.n40 PRE_CLSA.t1 718.909
R10045 PRE_CLSA.n38 PRE_CLSA.t97 718.909
R10046 PRE_CLSA.n36 PRE_CLSA.t25 718.909
R10047 PRE_CLSA.n34 PRE_CLSA.t91 718.909
R10048 PRE_CLSA.n32 PRE_CLSA.t122 718.909
R10049 PRE_CLSA.n31 PRE_CLSA.t59 718.909
R10050 PRE_CLSA.n94 PRE_CLSA.n30 30.983
R10051 PRE_CLSA.n126 PRE_CLSA.n94 24.254
R10052 PRE_CLSA.n33 PRE_CLSA.n31 16.71
R10053 PRE_CLSA.n93 PRE_CLSA.n92 13.414
R10054 PRE_CLSA.n91 PRE_CLSA.n90 13.414
R10055 PRE_CLSA.n89 PRE_CLSA.n88 13.414
R10056 PRE_CLSA.n87 PRE_CLSA.n86 13.414
R10057 PRE_CLSA.n85 PRE_CLSA.n84 13.414
R10058 PRE_CLSA.n83 PRE_CLSA.n82 13.414
R10059 PRE_CLSA.n81 PRE_CLSA.n80 13.414
R10060 PRE_CLSA.n79 PRE_CLSA.n78 13.414
R10061 PRE_CLSA.n77 PRE_CLSA.n76 13.414
R10062 PRE_CLSA.n75 PRE_CLSA.n74 13.414
R10063 PRE_CLSA.n73 PRE_CLSA.n72 13.414
R10064 PRE_CLSA.n71 PRE_CLSA.n70 13.414
R10065 PRE_CLSA.n69 PRE_CLSA.n68 13.414
R10066 PRE_CLSA.n67 PRE_CLSA.n66 13.414
R10067 PRE_CLSA.n65 PRE_CLSA.n64 13.414
R10068 PRE_CLSA.n63 PRE_CLSA.n62 13.414
R10069 PRE_CLSA.n61 PRE_CLSA.n60 13.414
R10070 PRE_CLSA.n59 PRE_CLSA.n58 13.414
R10071 PRE_CLSA.n57 PRE_CLSA.n56 13.414
R10072 PRE_CLSA.n55 PRE_CLSA.n54 13.414
R10073 PRE_CLSA.n53 PRE_CLSA.n52 13.414
R10074 PRE_CLSA.n51 PRE_CLSA.n50 13.414
R10075 PRE_CLSA.n49 PRE_CLSA.n48 13.414
R10076 PRE_CLSA.n47 PRE_CLSA.n46 13.414
R10077 PRE_CLSA.n45 PRE_CLSA.n44 13.414
R10078 PRE_CLSA.n43 PRE_CLSA.n42 13.414
R10079 PRE_CLSA.n41 PRE_CLSA.n40 13.414
R10080 PRE_CLSA.n39 PRE_CLSA.n38 13.414
R10081 PRE_CLSA.n37 PRE_CLSA.n36 13.414
R10082 PRE_CLSA.n35 PRE_CLSA.n34 13.414
R10083 PRE_CLSA.n33 PRE_CLSA.n32 13.414
R10084 PRE_CLSA.n98 PRE_CLSA.n97 6.883
R10085 PRE_CLSA.n100 PRE_CLSA.n99 6.883
R10086 PRE_CLSA.n3 PRE_CLSA.n2 6.883
R10087 PRE_CLSA.n5 PRE_CLSA.n4 6.883
R10088 PRE_CLSA.n102 PRE_CLSA.n101 6.856
R10089 PRE_CLSA.n104 PRE_CLSA.n103 6.856
R10090 PRE_CLSA.n7 PRE_CLSA.n6 6.856
R10091 PRE_CLSA.n9 PRE_CLSA.n8 6.856
R10092 PRE_CLSA.n106 PRE_CLSA.n105 6.838
R10093 PRE_CLSA.n108 PRE_CLSA.n107 6.838
R10094 PRE_CLSA.n110 PRE_CLSA.n109 6.838
R10095 PRE_CLSA.n112 PRE_CLSA.n111 6.838
R10096 PRE_CLSA.n114 PRE_CLSA.n113 6.838
R10097 PRE_CLSA.n116 PRE_CLSA.n115 6.838
R10098 PRE_CLSA.n122 PRE_CLSA.n121 6.838
R10099 PRE_CLSA.n11 PRE_CLSA.n10 6.838
R10100 PRE_CLSA.n13 PRE_CLSA.n12 6.838
R10101 PRE_CLSA.n15 PRE_CLSA.n14 6.838
R10102 PRE_CLSA.n17 PRE_CLSA.n16 6.838
R10103 PRE_CLSA.n19 PRE_CLSA.n18 6.838
R10104 PRE_CLSA.n21 PRE_CLSA.n20 6.838
R10105 PRE_CLSA.n27 PRE_CLSA.n26 6.838
R10106 PRE_CLSA.n118 PRE_CLSA.n117 6.829
R10107 PRE_CLSA.n120 PRE_CLSA.n119 6.829
R10108 PRE_CLSA.n23 PRE_CLSA.n22 6.829
R10109 PRE_CLSA.n25 PRE_CLSA.n24 6.829
R10110 PRE_CLSA.n126 PRE_CLSA.n125 6.724
R10111 PRE_CLSA.n94 PRE_CLSA.n93 6.579
R10112 PRE_CLSA.n124 PRE_CLSA.n123 6.553
R10113 PRE_CLSA.n29 PRE_CLSA.n28 6.553
R10114 PRE_CLSA.n39 PRE_CLSA.n37 6.437
R10115 PRE_CLSA.n43 PRE_CLSA.n41 6.437
R10116 PRE_CLSA.n47 PRE_CLSA.n45 6.412
R10117 PRE_CLSA.n51 PRE_CLSA.n49 6.412
R10118 PRE_CLSA.n55 PRE_CLSA.n53 6.396
R10119 PRE_CLSA.n59 PRE_CLSA.n57 6.396
R10120 PRE_CLSA.n63 PRE_CLSA.n61 6.396
R10121 PRE_CLSA.n67 PRE_CLSA.n65 6.396
R10122 PRE_CLSA.n71 PRE_CLSA.n69 6.396
R10123 PRE_CLSA.n75 PRE_CLSA.n73 6.396
R10124 PRE_CLSA.n87 PRE_CLSA.n85 6.396
R10125 PRE_CLSA.n79 PRE_CLSA.n77 6.387
R10126 PRE_CLSA.n83 PRE_CLSA.n81 6.387
R10127 PRE_CLSA.n91 PRE_CLSA.n89 6.129
R10128 PRE_CLSA.n96 PRE_CLSA.n95 4.329
R10129 PRE_CLSA.n1 PRE_CLSA.n0 4.329
R10130 PRE_CLSA.n35 PRE_CLSA.n33 4.054
R10131 PRE_CLSA PRE_CLSA.n126 3.678
R10132 PRE_CLSA.n97 PRE_CLSA.n96 3.517
R10133 PRE_CLSA.n99 PRE_CLSA.n98 3.517
R10134 PRE_CLSA.n101 PRE_CLSA.n100 3.517
R10135 PRE_CLSA.n103 PRE_CLSA.n102 3.517
R10136 PRE_CLSA.n105 PRE_CLSA.n104 3.517
R10137 PRE_CLSA.n107 PRE_CLSA.n106 3.517
R10138 PRE_CLSA.n109 PRE_CLSA.n108 3.517
R10139 PRE_CLSA.n111 PRE_CLSA.n110 3.517
R10140 PRE_CLSA.n113 PRE_CLSA.n112 3.517
R10141 PRE_CLSA.n115 PRE_CLSA.n114 3.517
R10142 PRE_CLSA.n117 PRE_CLSA.n116 3.517
R10143 PRE_CLSA.n119 PRE_CLSA.n118 3.517
R10144 PRE_CLSA.n121 PRE_CLSA.n120 3.517
R10145 PRE_CLSA.n123 PRE_CLSA.n122 3.517
R10146 PRE_CLSA.n125 PRE_CLSA.n124 3.517
R10147 PRE_CLSA.n2 PRE_CLSA.n1 3.517
R10148 PRE_CLSA.n4 PRE_CLSA.n3 3.517
R10149 PRE_CLSA.n6 PRE_CLSA.n5 3.517
R10150 PRE_CLSA.n8 PRE_CLSA.n7 3.517
R10151 PRE_CLSA.n10 PRE_CLSA.n9 3.517
R10152 PRE_CLSA.n12 PRE_CLSA.n11 3.517
R10153 PRE_CLSA.n14 PRE_CLSA.n13 3.517
R10154 PRE_CLSA.n16 PRE_CLSA.n15 3.517
R10155 PRE_CLSA.n18 PRE_CLSA.n17 3.517
R10156 PRE_CLSA.n20 PRE_CLSA.n19 3.517
R10157 PRE_CLSA.n22 PRE_CLSA.n21 3.517
R10158 PRE_CLSA.n24 PRE_CLSA.n23 3.517
R10159 PRE_CLSA.n26 PRE_CLSA.n25 3.517
R10160 PRE_CLSA.n28 PRE_CLSA.n27 3.517
R10161 PRE_CLSA.n30 PRE_CLSA.n29 3.517
R10162 PRE_CLSA.n37 PRE_CLSA.n35 3.296
R10163 PRE_CLSA.n41 PRE_CLSA.n39 3.296
R10164 PRE_CLSA.n45 PRE_CLSA.n43 3.296
R10165 PRE_CLSA.n49 PRE_CLSA.n47 3.296
R10166 PRE_CLSA.n53 PRE_CLSA.n51 3.296
R10167 PRE_CLSA.n57 PRE_CLSA.n55 3.296
R10168 PRE_CLSA.n61 PRE_CLSA.n59 3.296
R10169 PRE_CLSA.n65 PRE_CLSA.n63 3.296
R10170 PRE_CLSA.n69 PRE_CLSA.n67 3.296
R10171 PRE_CLSA.n73 PRE_CLSA.n71 3.296
R10172 PRE_CLSA.n77 PRE_CLSA.n75 3.296
R10173 PRE_CLSA.n81 PRE_CLSA.n79 3.296
R10174 PRE_CLSA.n85 PRE_CLSA.n83 3.296
R10175 PRE_CLSA.n89 PRE_CLSA.n87 3.296
R10176 PRE_CLSA.n93 PRE_CLSA.n91 3.296
R10177 a_n52_n8583.n0 a_n52_n8583.t4 1465.51
R10178 a_n52_n8583.n0 a_n52_n8583.t3 712.44
R10179 a_n52_n8583.n1 a_n52_n8583.t0 375.067
R10180 a_n52_n8583.n1 a_n52_n8583.t1 272.668
R10181 a_n52_n8583.n2 a_n52_n8583.n0 143.764
R10182 a_n52_n8583.t2 a_n52_n8583.n2 78.193
R10183 a_n52_n8583.n2 a_n52_n8583.n1 4.517
R10184 a_4972_n812.n0 a_4972_n812.t1 358.166
R10185 a_4972_n812.t4 a_4972_n812.t3 337.399
R10186 a_4972_n812.t3 a_4972_n812.t5 285.986
R10187 a_4972_n812.n0 a_4972_n812.t4 282.573
R10188 a_4972_n812.n1 a_4972_n812.t2 202.857
R10189 a_4972_n812.n1 a_4972_n812.n0 173.817
R10190 a_4972_n812.n1 a_4972_n812.t0 20.826
R10191 a_4972_n812.n2 a_4972_n812.n1 20.689
R10192 a_4877_n827.n0 a_4877_n827.t1 362.857
R10193 a_4877_n827.t4 a_4877_n827.t3 337.399
R10194 a_4877_n827.t3 a_4877_n827.t5 298.839
R10195 a_4877_n827.n0 a_4877_n827.t4 280.405
R10196 a_4877_n827.n1 a_4877_n827.t2 200
R10197 a_4877_n827.n1 a_4877_n827.n0 172.311
R10198 a_4877_n827.n2 a_4877_n827.n1 24
R10199 a_4877_n827.n1 a_4877_n827.t0 21.212
R10200 a_2590_n953.t35 a_2590_n953.n46 176.385
R10201 a_2590_n953.n22 a_2590_n953.t11 67.378
R10202 a_2590_n953.n0 a_2590_n953.t17 66.92
R10203 a_2590_n953.n1 a_2590_n953.t9 66.92
R10204 a_2590_n953.n2 a_2590_n953.t16 66.92
R10205 a_2590_n953.n3 a_2590_n953.t12 66.92
R10206 a_2590_n953.n4 a_2590_n953.t23 66.92
R10207 a_2590_n953.n5 a_2590_n953.t46 66.92
R10208 a_2590_n953.n6 a_2590_n953.t39 66.92
R10209 a_2590_n953.n7 a_2590_n953.t42 66.92
R10210 a_2590_n953.n8 a_2590_n953.t24 66.92
R10211 a_2590_n953.n9 a_2590_n953.t2 66.92
R10212 a_2590_n953.n10 a_2590_n953.t19 66.92
R10213 a_2590_n953.n11 a_2590_n953.t31 66.92
R10214 a_2590_n953.n12 a_2590_n953.t26 66.92
R10215 a_2590_n953.n13 a_2590_n953.t32 66.92
R10216 a_2590_n953.n14 a_2590_n953.t45 66.92
R10217 a_2590_n953.n15 a_2590_n953.t44 66.92
R10218 a_2590_n953.n16 a_2590_n953.t41 66.92
R10219 a_2590_n953.n17 a_2590_n953.t1 66.92
R10220 a_2590_n953.n18 a_2590_n953.t21 66.92
R10221 a_2590_n953.n19 a_2590_n953.t0 66.92
R10222 a_2590_n953.n20 a_2590_n953.t13 66.92
R10223 a_2590_n953.n21 a_2590_n953.t15 66.92
R10224 a_2590_n953.n22 a_2590_n953.t7 66.92
R10225 a_2590_n953.n23 a_2590_n953.t14 65.518
R10226 a_2590_n953.n45 a_2590_n953.t18 63.519
R10227 a_2590_n953.n44 a_2590_n953.t5 63.519
R10228 a_2590_n953.n43 a_2590_n953.t10 63.519
R10229 a_2590_n953.n42 a_2590_n953.t3 63.519
R10230 a_2590_n953.n41 a_2590_n953.t30 63.519
R10231 a_2590_n953.n40 a_2590_n953.t38 63.519
R10232 a_2590_n953.n39 a_2590_n953.t22 63.519
R10233 a_2590_n953.n38 a_2590_n953.t20 63.519
R10234 a_2590_n953.n37 a_2590_n953.t43 63.519
R10235 a_2590_n953.n36 a_2590_n953.t37 63.519
R10236 a_2590_n953.n35 a_2590_n953.t29 63.519
R10237 a_2590_n953.n34 a_2590_n953.t28 63.519
R10238 a_2590_n953.n33 a_2590_n953.t33 63.519
R10239 a_2590_n953.n32 a_2590_n953.t40 63.519
R10240 a_2590_n953.n31 a_2590_n953.t47 63.519
R10241 a_2590_n953.n30 a_2590_n953.t36 63.519
R10242 a_2590_n953.n29 a_2590_n953.t34 63.519
R10243 a_2590_n953.n28 a_2590_n953.t48 63.519
R10244 a_2590_n953.n27 a_2590_n953.t27 63.519
R10245 a_2590_n953.n26 a_2590_n953.t25 63.519
R10246 a_2590_n953.n25 a_2590_n953.t8 63.519
R10247 a_2590_n953.n24 a_2590_n953.t6 63.519
R10248 a_2590_n953.n23 a_2590_n953.t4 63.519
R10249 a_2590_n953.n46 a_2590_n953.n0 19.599
R10250 a_2590_n953.n46 a_2590_n953.n45 15.67
R10251 a_2590_n953.n44 a_2590_n953.n43 2.524
R10252 a_2590_n953.n24 a_2590_n953.n23 2.498
R10253 a_2590_n953.n21 a_2590_n953.n22 2.495
R10254 a_2590_n953.n1 a_2590_n953.n2 2.459
R10255 a_2590_n953.n38 a_2590_n953.n37 2.364
R10256 a_2590_n953.n30 a_2590_n953.n29 2.355
R10257 a_2590_n953.n7 a_2590_n953.n8 2.299
R10258 a_2590_n953.n15 a_2590_n953.n16 2.29
R10259 a_2590_n953.n16 a_2590_n953.n17 2.057
R10260 a_2590_n953.n8 a_2590_n953.n9 2.057
R10261 a_2590_n953.n2 a_2590_n953.n3 2.057
R10262 a_2590_n953.n0 a_2590_n953.n1 2.057
R10263 a_2590_n953.n45 a_2590_n953.n44 1.998
R10264 a_2590_n953.n43 a_2590_n953.n42 1.998
R10265 a_2590_n953.n42 a_2590_n953.n41 1.998
R10266 a_2590_n953.n41 a_2590_n953.n40 1.998
R10267 a_2590_n953.n40 a_2590_n953.n39 1.998
R10268 a_2590_n953.n39 a_2590_n953.n38 1.998
R10269 a_2590_n953.n37 a_2590_n953.n36 1.998
R10270 a_2590_n953.n36 a_2590_n953.n35 1.998
R10271 a_2590_n953.n35 a_2590_n953.n34 1.998
R10272 a_2590_n953.n34 a_2590_n953.n33 1.998
R10273 a_2590_n953.n33 a_2590_n953.n32 1.998
R10274 a_2590_n953.n32 a_2590_n953.n31 1.998
R10275 a_2590_n953.n31 a_2590_n953.n30 1.998
R10276 a_2590_n953.n29 a_2590_n953.n28 1.998
R10277 a_2590_n953.n28 a_2590_n953.n27 1.998
R10278 a_2590_n953.n27 a_2590_n953.n26 1.998
R10279 a_2590_n953.n26 a_2590_n953.n25 1.998
R10280 a_2590_n953.n25 a_2590_n953.n24 1.998
R10281 a_2590_n953.n20 a_2590_n953.n21 1.995
R10282 a_2590_n953.n19 a_2590_n953.n20 1.995
R10283 a_2590_n953.n18 a_2590_n953.n19 1.995
R10284 a_2590_n953.n17 a_2590_n953.n18 1.995
R10285 a_2590_n953.n14 a_2590_n953.n15 1.995
R10286 a_2590_n953.n13 a_2590_n953.n14 1.995
R10287 a_2590_n953.n12 a_2590_n953.n13 1.995
R10288 a_2590_n953.n11 a_2590_n953.n12 1.995
R10289 a_2590_n953.n10 a_2590_n953.n11 1.995
R10290 a_2590_n953.n9 a_2590_n953.n10 1.995
R10291 a_2590_n953.n6 a_2590_n953.n7 1.995
R10292 a_2590_n953.n5 a_2590_n953.n6 1.995
R10293 a_2590_n953.n4 a_2590_n953.n5 1.995
R10294 a_2590_n953.n3 a_2590_n953.n4 1.995
R10295 a_3042_4445.t0 a_3042_4445.t1 242.857
R10296 a_5452_196.n0 a_5452_196.t1 362.857
R10297 a_5452_196.t3 a_5452_196.t5 337.399
R10298 a_5452_196.t5 a_5452_196.t4 298.839
R10299 a_5452_196.n0 a_5452_196.t3 280.405
R10300 a_5452_196.n1 a_5452_196.t2 200
R10301 a_5452_196.n1 a_5452_196.n0 172.311
R10302 a_5452_196.n2 a_5452_196.n1 24
R10303 a_5452_196.n1 a_5452_196.t0 21.212
R10304 a_5547_211.n0 a_5547_211.t1 358.166
R10305 a_5547_211.t4 a_5547_211.t3 337.399
R10306 a_5547_211.t3 a_5547_211.t5 285.986
R10307 a_5547_211.n0 a_5547_211.t4 282.573
R10308 a_5547_211.n1 a_5547_211.t2 202.857
R10309 a_5547_211.n1 a_5547_211.n0 173.817
R10310 a_5547_211.n1 a_5547_211.t0 20.826
R10311 a_5547_211.n2 a_5547_211.n1 20.689
R10312 a_2672_n30.n0 a_2672_n30.t0 358.166
R10313 a_2672_n30.t3 a_2672_n30.t4 337.399
R10314 a_2672_n30.t4 a_2672_n30.t5 285.986
R10315 a_2672_n30.n0 a_2672_n30.t3 282.573
R10316 a_2672_n30.n1 a_2672_n30.t2 202.857
R10317 a_2672_n30.n1 a_2672_n30.n0 173.817
R10318 a_2672_n30.n1 a_2672_n30.t1 20.826
R10319 a_2672_n30.n2 a_2672_n30.n1 20.689
R10320 a_2577_n45.n0 a_2577_n45.t1 362.857
R10321 a_2577_n45.t5 a_2577_n45.t4 337.399
R10322 a_2577_n45.t4 a_2577_n45.t3 298.839
R10323 a_2577_n45.n0 a_2577_n45.t5 280.405
R10324 a_2577_n45.n1 a_2577_n45.t2 200
R10325 a_2577_n45.n1 a_2577_n45.n0 172.311
R10326 a_2577_n45.n2 a_2577_n45.n1 24
R10327 a_2577_n45.n1 a_2577_n45.t0 21.212
R10328 a_6697_n271.n0 a_6697_n271.t0 358.166
R10329 a_6697_n271.t5 a_6697_n271.t3 337.399
R10330 a_6697_n271.t3 a_6697_n271.t4 285.986
R10331 a_6697_n271.n0 a_6697_n271.t5 282.573
R10332 a_6697_n271.n1 a_6697_n271.t2 202.857
R10333 a_6697_n271.n1 a_6697_n271.n0 173.817
R10334 a_6697_n271.n1 a_6697_n271.t1 20.826
R10335 a_6697_n271.n2 a_6697_n271.n1 20.689
R10336 a_6602_n286.n0 a_6602_n286.t1 362.857
R10337 a_6602_n286.t3 a_6602_n286.t5 337.399
R10338 a_6602_n286.t5 a_6602_n286.t4 298.839
R10339 a_6602_n286.n0 a_6602_n286.t3 280.405
R10340 a_6602_n286.n1 a_6602_n286.t2 200
R10341 a_6602_n286.n1 a_6602_n286.n0 172.311
R10342 a_6602_n286.n2 a_6602_n286.n1 24
R10343 a_6602_n286.n1 a_6602_n286.t0 21.212
R10344 a_4315_4445.t0 a_4315_4445.t1 242.857
R10345 a_4315_n953.t32 a_4315_n953.n46 176.385
R10346 a_4315_n953.n22 a_4315_n953.t11 67.378
R10347 a_4315_n953.n0 a_4315_n953.t17 66.92
R10348 a_4315_n953.n1 a_4315_n953.t3 66.92
R10349 a_4315_n953.n2 a_4315_n953.t8 66.92
R10350 a_4315_n953.n3 a_4315_n953.t16 66.92
R10351 a_4315_n953.n4 a_4315_n953.t2 66.92
R10352 a_4315_n953.n5 a_4315_n953.t1 66.92
R10353 a_4315_n953.n6 a_4315_n953.t37 66.92
R10354 a_4315_n953.n7 a_4315_n953.t39 66.92
R10355 a_4315_n953.n8 a_4315_n953.t23 66.92
R10356 a_4315_n953.n9 a_4315_n953.t0 66.92
R10357 a_4315_n953.n10 a_4315_n953.t19 66.92
R10358 a_4315_n953.n11 a_4315_n953.t30 66.92
R10359 a_4315_n953.n12 a_4315_n953.t25 66.92
R10360 a_4315_n953.n13 a_4315_n953.t41 66.92
R10361 a_4315_n953.n14 a_4315_n953.t48 66.92
R10362 a_4315_n953.n15 a_4315_n953.t44 66.92
R10363 a_4315_n953.n16 a_4315_n953.t45 66.92
R10364 a_4315_n953.n17 a_4315_n953.t46 66.92
R10365 a_4315_n953.n18 a_4315_n953.t21 66.92
R10366 a_4315_n953.n19 a_4315_n953.t47 66.92
R10367 a_4315_n953.n20 a_4315_n953.t12 66.92
R10368 a_4315_n953.n21 a_4315_n953.t7 66.92
R10369 a_4315_n953.n22 a_4315_n953.t5 66.92
R10370 a_4315_n953.n23 a_4315_n953.t10 65.518
R10371 a_4315_n953.n45 a_4315_n953.t4 63.519
R10372 a_4315_n953.n44 a_4315_n953.t15 63.519
R10373 a_4315_n953.n43 a_4315_n953.t13 63.519
R10374 a_4315_n953.n42 a_4315_n953.t6 63.519
R10375 a_4315_n953.n41 a_4315_n953.t29 63.519
R10376 a_4315_n953.n40 a_4315_n953.t36 63.519
R10377 a_4315_n953.n39 a_4315_n953.t22 63.519
R10378 a_4315_n953.n38 a_4315_n953.t20 63.519
R10379 a_4315_n953.n37 a_4315_n953.t43 63.519
R10380 a_4315_n953.n36 a_4315_n953.t35 63.519
R10381 a_4315_n953.n35 a_4315_n953.t28 63.519
R10382 a_4315_n953.n34 a_4315_n953.t27 63.519
R10383 a_4315_n953.n33 a_4315_n953.t33 63.519
R10384 a_4315_n953.n32 a_4315_n953.t38 63.519
R10385 a_4315_n953.n31 a_4315_n953.t40 63.519
R10386 a_4315_n953.n30 a_4315_n953.t34 63.519
R10387 a_4315_n953.n29 a_4315_n953.t31 63.519
R10388 a_4315_n953.n28 a_4315_n953.t42 63.519
R10389 a_4315_n953.n27 a_4315_n953.t26 63.519
R10390 a_4315_n953.n26 a_4315_n953.t24 63.519
R10391 a_4315_n953.n25 a_4315_n953.t9 63.519
R10392 a_4315_n953.n24 a_4315_n953.t14 63.519
R10393 a_4315_n953.n23 a_4315_n953.t18 63.519
R10394 a_4315_n953.n46 a_4315_n953.n45 18.144
R10395 a_4315_n953.n46 a_4315_n953.n0 17.125
R10396 a_4315_n953.n44 a_4315_n953.n43 2.524
R10397 a_4315_n953.n24 a_4315_n953.n23 2.498
R10398 a_4315_n953.n21 a_4315_n953.n22 2.495
R10399 a_4315_n953.n1 a_4315_n953.n2 2.459
R10400 a_4315_n953.n38 a_4315_n953.n37 2.364
R10401 a_4315_n953.n30 a_4315_n953.n29 2.355
R10402 a_4315_n953.n7 a_4315_n953.n8 2.299
R10403 a_4315_n953.n15 a_4315_n953.n16 2.29
R10404 a_4315_n953.n16 a_4315_n953.n17 2.057
R10405 a_4315_n953.n8 a_4315_n953.n9 2.057
R10406 a_4315_n953.n2 a_4315_n953.n3 2.057
R10407 a_4315_n953.n0 a_4315_n953.n1 2.057
R10408 a_4315_n953.n45 a_4315_n953.n44 1.998
R10409 a_4315_n953.n43 a_4315_n953.n42 1.998
R10410 a_4315_n953.n42 a_4315_n953.n41 1.998
R10411 a_4315_n953.n41 a_4315_n953.n40 1.998
R10412 a_4315_n953.n40 a_4315_n953.n39 1.998
R10413 a_4315_n953.n39 a_4315_n953.n38 1.998
R10414 a_4315_n953.n37 a_4315_n953.n36 1.998
R10415 a_4315_n953.n36 a_4315_n953.n35 1.998
R10416 a_4315_n953.n35 a_4315_n953.n34 1.998
R10417 a_4315_n953.n34 a_4315_n953.n33 1.998
R10418 a_4315_n953.n33 a_4315_n953.n32 1.998
R10419 a_4315_n953.n32 a_4315_n953.n31 1.998
R10420 a_4315_n953.n31 a_4315_n953.n30 1.998
R10421 a_4315_n953.n29 a_4315_n953.n28 1.998
R10422 a_4315_n953.n28 a_4315_n953.n27 1.998
R10423 a_4315_n953.n27 a_4315_n953.n26 1.998
R10424 a_4315_n953.n26 a_4315_n953.n25 1.998
R10425 a_4315_n953.n25 a_4315_n953.n24 1.998
R10426 a_4315_n953.n20 a_4315_n953.n21 1.995
R10427 a_4315_n953.n19 a_4315_n953.n20 1.995
R10428 a_4315_n953.n18 a_4315_n953.n19 1.995
R10429 a_4315_n953.n17 a_4315_n953.n18 1.995
R10430 a_4315_n953.n14 a_4315_n953.n15 1.995
R10431 a_4315_n953.n13 a_4315_n953.n14 1.995
R10432 a_4315_n953.n12 a_4315_n953.n13 1.995
R10433 a_4315_n953.n11 a_4315_n953.n12 1.995
R10434 a_4315_n953.n10 a_4315_n953.n11 1.995
R10435 a_4315_n953.n9 a_4315_n953.n10 1.995
R10436 a_4315_n953.n6 a_4315_n953.n7 1.995
R10437 a_4315_n953.n5 a_4315_n953.n6 1.995
R10438 a_4315_n953.n4 a_4315_n953.n5 1.995
R10439 a_4315_n953.n3 a_4315_n953.n4 1.995
R10440 SA_OUT[10].n1 SA_OUT[10].t4 661.027
R10441 SA_OUT[10].n1 SA_OUT[10].t3 392.255
R10442 SA_OUT[10].n2 SA_OUT[10].t0 223.716
R10443 SA_OUT[10].n0 SA_OUT[10].t2 153.977
R10444 SA_OUT[10].n2 SA_OUT[10].n1 143.764
R10445 SA_OUT[10].n0 SA_OUT[10].t1 59.86
R10446 SA_OUT[10] SA_OUT[10].n3 14.537
R10447 SA_OUT[10].n3 SA_OUT[10].n0 3.011
R10448 SA_OUT[10].n3 SA_OUT[10].n2 1.505
R10449 a_7190_n512.t0 a_7190_n512.t1 242.857
R10450 a_7190_n953.t32 a_7190_n953.n46 176.385
R10451 a_7190_n953.n22 a_7190_n953.t9 67.378
R10452 a_7190_n953.n0 a_7190_n953.t11 66.92
R10453 a_7190_n953.n1 a_7190_n953.t18 66.92
R10454 a_7190_n953.n2 a_7190_n953.t7 66.92
R10455 a_7190_n953.n3 a_7190_n953.t4 66.92
R10456 a_7190_n953.n4 a_7190_n953.t3 66.92
R10457 a_7190_n953.n5 a_7190_n953.t48 66.92
R10458 a_7190_n953.n6 a_7190_n953.t38 66.92
R10459 a_7190_n953.n7 a_7190_n953.t42 66.92
R10460 a_7190_n953.n8 a_7190_n953.t24 66.92
R10461 a_7190_n953.n9 a_7190_n953.t2 66.92
R10462 a_7190_n953.n10 a_7190_n953.t20 66.92
R10463 a_7190_n953.n11 a_7190_n953.t29 66.92
R10464 a_7190_n953.n12 a_7190_n953.t26 66.92
R10465 a_7190_n953.n13 a_7190_n953.t44 66.92
R10466 a_7190_n953.n14 a_7190_n953.t47 66.92
R10467 a_7190_n953.n15 a_7190_n953.t46 66.92
R10468 a_7190_n953.n16 a_7190_n953.t40 66.92
R10469 a_7190_n953.n17 a_7190_n953.t0 66.92
R10470 a_7190_n953.n18 a_7190_n953.t23 66.92
R10471 a_7190_n953.n19 a_7190_n953.t1 66.92
R10472 a_7190_n953.n20 a_7190_n953.t8 66.92
R10473 a_7190_n953.n21 a_7190_n953.t14 66.92
R10474 a_7190_n953.n22 a_7190_n953.t17 66.92
R10475 a_7190_n953.n23 a_7190_n953.t12 65.518
R10476 a_7190_n953.n45 a_7190_n953.t10 63.519
R10477 a_7190_n953.n44 a_7190_n953.t16 63.519
R10478 a_7190_n953.n43 a_7190_n953.t13 63.519
R10479 a_7190_n953.n42 a_7190_n953.t19 63.519
R10480 a_7190_n953.n41 a_7190_n953.t33 63.519
R10481 a_7190_n953.n40 a_7190_n953.t37 63.519
R10482 a_7190_n953.n39 a_7190_n953.t22 63.519
R10483 a_7190_n953.n38 a_7190_n953.t21 63.519
R10484 a_7190_n953.n37 a_7190_n953.t41 63.519
R10485 a_7190_n953.n36 a_7190_n953.t36 63.519
R10486 a_7190_n953.n35 a_7190_n953.t28 63.519
R10487 a_7190_n953.n34 a_7190_n953.t30 63.519
R10488 a_7190_n953.n33 a_7190_n953.t34 63.519
R10489 a_7190_n953.n32 a_7190_n953.t39 63.519
R10490 a_7190_n953.n31 a_7190_n953.t43 63.519
R10491 a_7190_n953.n30 a_7190_n953.t35 63.519
R10492 a_7190_n953.n29 a_7190_n953.t31 63.519
R10493 a_7190_n953.n28 a_7190_n953.t45 63.519
R10494 a_7190_n953.n27 a_7190_n953.t27 63.519
R10495 a_7190_n953.n26 a_7190_n953.t25 63.519
R10496 a_7190_n953.n25 a_7190_n953.t15 63.519
R10497 a_7190_n953.n24 a_7190_n953.t6 63.519
R10498 a_7190_n953.n23 a_7190_n953.t5 63.519
R10499 a_7190_n953.n46 a_7190_n953.n0 19.599
R10500 a_7190_n953.n46 a_7190_n953.n45 15.67
R10501 a_7190_n953.n44 a_7190_n953.n43 2.524
R10502 a_7190_n953.n24 a_7190_n953.n23 2.498
R10503 a_7190_n953.n21 a_7190_n953.n22 2.495
R10504 a_7190_n953.n1 a_7190_n953.n2 2.459
R10505 a_7190_n953.n38 a_7190_n953.n37 2.364
R10506 a_7190_n953.n30 a_7190_n953.n29 2.355
R10507 a_7190_n953.n7 a_7190_n953.n8 2.299
R10508 a_7190_n953.n15 a_7190_n953.n16 2.29
R10509 a_7190_n953.n16 a_7190_n953.n17 2.057
R10510 a_7190_n953.n8 a_7190_n953.n9 2.057
R10511 a_7190_n953.n2 a_7190_n953.n3 2.057
R10512 a_7190_n953.n0 a_7190_n953.n1 2.057
R10513 a_7190_n953.n45 a_7190_n953.n44 1.998
R10514 a_7190_n953.n43 a_7190_n953.n42 1.998
R10515 a_7190_n953.n42 a_7190_n953.n41 1.998
R10516 a_7190_n953.n41 a_7190_n953.n40 1.998
R10517 a_7190_n953.n40 a_7190_n953.n39 1.998
R10518 a_7190_n953.n39 a_7190_n953.n38 1.998
R10519 a_7190_n953.n37 a_7190_n953.n36 1.998
R10520 a_7190_n953.n36 a_7190_n953.n35 1.998
R10521 a_7190_n953.n35 a_7190_n953.n34 1.998
R10522 a_7190_n953.n34 a_7190_n953.n33 1.998
R10523 a_7190_n953.n33 a_7190_n953.n32 1.998
R10524 a_7190_n953.n32 a_7190_n953.n31 1.998
R10525 a_7190_n953.n31 a_7190_n953.n30 1.998
R10526 a_7190_n953.n29 a_7190_n953.n28 1.998
R10527 a_7190_n953.n28 a_7190_n953.n27 1.998
R10528 a_7190_n953.n27 a_7190_n953.n26 1.998
R10529 a_7190_n953.n26 a_7190_n953.n25 1.998
R10530 a_7190_n953.n25 a_7190_n953.n24 1.998
R10531 a_7190_n953.n20 a_7190_n953.n21 1.995
R10532 a_7190_n953.n19 a_7190_n953.n20 1.995
R10533 a_7190_n953.n18 a_7190_n953.n19 1.995
R10534 a_7190_n953.n17 a_7190_n953.n18 1.995
R10535 a_7190_n953.n14 a_7190_n953.n15 1.995
R10536 a_7190_n953.n13 a_7190_n953.n14 1.995
R10537 a_7190_n953.n12 a_7190_n953.n13 1.995
R10538 a_7190_n953.n11 a_7190_n953.n12 1.995
R10539 a_7190_n953.n10 a_7190_n953.n11 1.995
R10540 a_7190_n953.n9 a_7190_n953.n10 1.995
R10541 a_7190_n953.n6 a_7190_n953.n7 1.995
R10542 a_7190_n953.n5 a_7190_n953.n6 1.995
R10543 a_7190_n953.n4 a_7190_n953.n5 1.995
R10544 a_7190_n953.n3 a_7190_n953.n4 1.995
R10545 WWL[10].n0 WWL[10].t15 262.032
R10546 WWL[10].n29 WWL[10].t18 260.715
R10547 WWL[10].n27 WWL[10].t21 260.715
R10548 WWL[10].n25 WWL[10].t3 260.715
R10549 WWL[10].n23 WWL[10].t29 260.715
R10550 WWL[10].n21 WWL[10].t9 260.715
R10551 WWL[10].n19 WWL[10].t26 260.715
R10552 WWL[10].n17 WWL[10].t17 260.715
R10553 WWL[10].n15 WWL[10].t0 260.715
R10554 WWL[10].n13 WWL[10].t22 260.715
R10555 WWL[10].n11 WWL[10].t30 260.715
R10556 WWL[10].n9 WWL[10].t19 260.715
R10557 WWL[10].n7 WWL[10].t1 260.715
R10558 WWL[10].n5 WWL[10].t27 260.715
R10559 WWL[10].n3 WWL[10].t10 260.715
R10560 WWL[10].n1 WWL[10].t23 260.715
R10561 WWL[10].n30 WWL[10].t2 259.254
R10562 WWL[10].n28 WWL[10].t8 259.254
R10563 WWL[10].n26 WWL[10].t20 259.254
R10564 WWL[10].n24 WWL[10].t4 259.254
R10565 WWL[10].n22 WWL[10].t28 259.254
R10566 WWL[10].n20 WWL[10].t11 259.254
R10567 WWL[10].n18 WWL[10].t24 259.254
R10568 WWL[10].n16 WWL[10].t6 259.254
R10569 WWL[10].n14 WWL[10].t31 259.254
R10570 WWL[10].n12 WWL[10].t14 259.254
R10571 WWL[10].n10 WWL[10].t5 259.254
R10572 WWL[10].n8 WWL[10].t12 259.254
R10573 WWL[10].n6 WWL[10].t13 259.254
R10574 WWL[10].n4 WWL[10].t16 259.254
R10575 WWL[10].n2 WWL[10].t7 259.254
R10576 WWL[10].n0 WWL[10].t25 259.254
R10577 WWL[10] WWL[10].n30 44.647
R10578 WWL[10].n1 WWL[10].n0 3.576
R10579 WWL[10].n3 WWL[10].n2 3.576
R10580 WWL[10].n5 WWL[10].n4 3.576
R10581 WWL[10].n7 WWL[10].n6 3.576
R10582 WWL[10].n9 WWL[10].n8 3.576
R10583 WWL[10].n11 WWL[10].n10 3.576
R10584 WWL[10].n13 WWL[10].n12 3.576
R10585 WWL[10].n15 WWL[10].n14 3.576
R10586 WWL[10].n17 WWL[10].n16 3.576
R10587 WWL[10].n19 WWL[10].n18 3.576
R10588 WWL[10].n21 WWL[10].n20 3.576
R10589 WWL[10].n23 WWL[10].n22 3.576
R10590 WWL[10].n25 WWL[10].n24 3.576
R10591 WWL[10].n27 WWL[10].n26 3.576
R10592 WWL[10].n29 WWL[10].n28 3.576
R10593 WWL[10].n2 WWL[10].n1 1.317
R10594 WWL[10].n4 WWL[10].n3 1.317
R10595 WWL[10].n6 WWL[10].n5 1.317
R10596 WWL[10].n8 WWL[10].n7 1.317
R10597 WWL[10].n10 WWL[10].n9 1.317
R10598 WWL[10].n12 WWL[10].n11 1.317
R10599 WWL[10].n14 WWL[10].n13 1.317
R10600 WWL[10].n16 WWL[10].n15 1.317
R10601 WWL[10].n18 WWL[10].n17 1.317
R10602 WWL[10].n20 WWL[10].n19 1.317
R10603 WWL[10].n22 WWL[10].n21 1.317
R10604 WWL[10].n24 WWL[10].n23 1.317
R10605 WWL[10].n26 WWL[10].n25 1.317
R10606 WWL[10].n28 WWL[10].n27 1.317
R10607 WWL[10].n30 WWL[10].n29 1.317
R10608 a_4570_4887.n25 a_4570_4887.t27 561.971
R10609 a_4570_4887.n0 a_4570_4887.t20 449.944
R10610 a_4570_4887.t24 a_4570_4887.n25 108.636
R10611 a_4570_4887.n0 a_4570_4887.t21 74.821
R10612 a_4570_4887.n24 a_4570_4887.t25 63.519
R10613 a_4570_4887.n23 a_4570_4887.t7 63.519
R10614 a_4570_4887.n22 a_4570_4887.t5 63.519
R10615 a_4570_4887.n21 a_4570_4887.t16 63.519
R10616 a_4570_4887.n20 a_4570_4887.t11 63.519
R10617 a_4570_4887.n19 a_4570_4887.t17 63.519
R10618 a_4570_4887.n18 a_4570_4887.t19 63.519
R10619 a_4570_4887.n17 a_4570_4887.t14 63.519
R10620 a_4570_4887.n16 a_4570_4887.t26 63.519
R10621 a_4570_4887.n15 a_4570_4887.t6 63.519
R10622 a_4570_4887.n14 a_4570_4887.t13 63.519
R10623 a_4570_4887.n13 a_4570_4887.t2 63.519
R10624 a_4570_4887.n12 a_4570_4887.t1 63.519
R10625 a_4570_4887.n11 a_4570_4887.t12 63.519
R10626 a_4570_4887.n10 a_4570_4887.t4 63.519
R10627 a_4570_4887.n9 a_4570_4887.t9 63.519
R10628 a_4570_4887.n8 a_4570_4887.t8 63.519
R10629 a_4570_4887.n7 a_4570_4887.t22 63.519
R10630 a_4570_4887.n6 a_4570_4887.t3 63.519
R10631 a_4570_4887.n5 a_4570_4887.t23 63.519
R10632 a_4570_4887.n4 a_4570_4887.t0 63.519
R10633 a_4570_4887.n3 a_4570_4887.t10 63.519
R10634 a_4570_4887.n2 a_4570_4887.t15 63.519
R10635 a_4570_4887.n1 a_4570_4887.t18 63.519
R10636 a_4570_4887.n1 a_4570_4887.n0 8.619
R10637 a_4570_4887.n25 a_4570_4887.n24 2.946
R10638 a_4570_4887.n23 a_4570_4887.n22 2.524
R10639 a_4570_4887.n3 a_4570_4887.n2 2.498
R10640 a_4570_4887.n17 a_4570_4887.n16 2.364
R10641 a_4570_4887.n9 a_4570_4887.n8 2.355
R10642 a_4570_4887.n24 a_4570_4887.n23 1.998
R10643 a_4570_4887.n22 a_4570_4887.n21 1.998
R10644 a_4570_4887.n21 a_4570_4887.n20 1.998
R10645 a_4570_4887.n20 a_4570_4887.n19 1.998
R10646 a_4570_4887.n19 a_4570_4887.n18 1.998
R10647 a_4570_4887.n18 a_4570_4887.n17 1.998
R10648 a_4570_4887.n16 a_4570_4887.n15 1.998
R10649 a_4570_4887.n15 a_4570_4887.n14 1.998
R10650 a_4570_4887.n14 a_4570_4887.n13 1.998
R10651 a_4570_4887.n13 a_4570_4887.n12 1.998
R10652 a_4570_4887.n12 a_4570_4887.n11 1.998
R10653 a_4570_4887.n11 a_4570_4887.n10 1.998
R10654 a_4570_4887.n10 a_4570_4887.n9 1.998
R10655 a_4570_4887.n8 a_4570_4887.n7 1.998
R10656 a_4570_4887.n7 a_4570_4887.n6 1.998
R10657 a_4570_4887.n6 a_4570_4887.n5 1.998
R10658 a_4570_4887.n5 a_4570_4887.n4 1.998
R10659 a_4570_4887.n4 a_4570_4887.n3 1.998
R10660 a_4570_4887.n2 a_4570_4887.n1 1.998
R10661 a_4302_1201.n0 a_4302_1201.t1 362.857
R10662 a_4302_1201.t3 a_4302_1201.t5 337.399
R10663 a_4302_1201.t5 a_4302_1201.t4 298.839
R10664 a_4302_1201.n0 a_4302_1201.t3 280.405
R10665 a_4302_1201.n1 a_4302_1201.t0 200
R10666 a_4302_1201.n1 a_4302_1201.n0 172.311
R10667 a_4302_1201.n2 a_4302_1201.n1 24
R10668 a_4302_1201.n1 a_4302_1201.t2 21.212
R10669 a_6602_960.n0 a_6602_960.t0 362.857
R10670 a_6602_960.t5 a_6602_960.t4 337.399
R10671 a_6602_960.t4 a_6602_960.t3 298.839
R10672 a_6602_960.n0 a_6602_960.t5 280.405
R10673 a_6602_960.n1 a_6602_960.t2 200
R10674 a_6602_960.n1 a_6602_960.n0 172.311
R10675 a_6602_960.n2 a_6602_960.n1 24
R10676 a_6602_960.n1 a_6602_960.t1 21.212
R10677 a_6615_975.t0 a_6615_975.t1 242.857
R10678 a_n3827_n4378.n3 a_n3827_n4378.t2 476.143
R10679 a_n3827_n4378.t6 a_n3827_n4378.t4 228.696
R10680 a_n3827_n4378.n2 a_n3827_n4378.t1 185.704
R10681 a_n3827_n4378.n0 a_n3827_n4378.t6 126.761
R10682 a_n3827_n4378.n1 a_n3827_n4378.t7 126.284
R10683 a_n3827_n4378.n1 a_n3827_n4378.t0 126.284
R10684 a_n3827_n4378.t3 a_n3827_n4378.n3 124.375
R10685 a_n3827_n4378.t0 a_n3827_n4378.n0 115.122
R10686 a_n3827_n4378.n3 a_n3827_n4378.n2 114.784
R10687 a_n3827_n4378.n0 a_n3827_n4378.t5 111.229
R10688 a_n3827_n4378.n2 a_n3827_n4378.n1 8.764
R10689 a_n3827_n7825.t0 a_n3827_n7825.t1 42.705
R10690 VCLP.n79 VCLP.t56 1367.97
R10691 VCLP.n31 VCLP.t36 1367.97
R10692 VCLP.n63 VCLP.t58 1366.51
R10693 VCLP.n0 VCLP.t92 1366.51
R10694 VCLP.n108 VCLP.t89 1365.35
R10695 VCLP.n106 VCLP.t13 1365.35
R10696 VCLP.n104 VCLP.t77 1365.35
R10697 VCLP.n102 VCLP.t78 1365.35
R10698 VCLP.n100 VCLP.t66 1365.35
R10699 VCLP.n98 VCLP.t27 1365.35
R10700 VCLP.n96 VCLP.t70 1365.35
R10701 VCLP.n94 VCLP.t31 1365.35
R10702 VCLP.n92 VCLP.t72 1365.35
R10703 VCLP.n90 VCLP.t34 1365.35
R10704 VCLP.n88 VCLP.t110 1365.35
R10705 VCLP.n86 VCLP.t81 1365.35
R10706 VCLP.n84 VCLP.t85 1365.35
R10707 VCLP.n82 VCLP.t106 1365.35
R10708 VCLP.n80 VCLP.t88 1365.35
R10709 VCLP.n60 VCLP.t63 1365.35
R10710 VCLP.n58 VCLP.t102 1365.35
R10711 VCLP.n56 VCLP.t50 1365.35
R10712 VCLP.n54 VCLP.t51 1365.35
R10713 VCLP.n52 VCLP.t40 1365.35
R10714 VCLP.n50 VCLP.t8 1365.35
R10715 VCLP.n48 VCLP.t45 1365.35
R10716 VCLP.n46 VCLP.t10 1365.35
R10717 VCLP.n44 VCLP.t46 1365.35
R10718 VCLP.n42 VCLP.t11 1365.35
R10719 VCLP.n40 VCLP.t87 1365.35
R10720 VCLP.n38 VCLP.t54 1365.35
R10721 VCLP.n36 VCLP.t59 1365.35
R10722 VCLP.n34 VCLP.t82 1365.35
R10723 VCLP.n32 VCLP.t60 1365.35
R10724 VCLP.n76 VCLP.t3 1363.89
R10725 VCLP.n74 VCLP.t39 1363.89
R10726 VCLP.n72 VCLP.t103 1363.89
R10727 VCLP.n70 VCLP.t104 1363.89
R10728 VCLP.n68 VCLP.t94 1363.89
R10729 VCLP.n66 VCLP.t55 1363.89
R10730 VCLP.n64 VCLP.t97 1363.89
R10731 VCLP.n29 VCLP.t7 1363.89
R10732 VCLP.n27 VCLP.t43 1363.89
R10733 VCLP.n25 VCLP.t108 1363.89
R10734 VCLP.n23 VCLP.t109 1363.89
R10735 VCLP.n21 VCLP.t96 1363.89
R10736 VCLP.n19 VCLP.t57 1363.89
R10737 VCLP.n17 VCLP.t100 1363.89
R10738 VCLP.n15 VCLP.t62 1363.89
R10739 VCLP.n13 VCLP.t101 1363.89
R10740 VCLP.n11 VCLP.t64 1363.89
R10741 VCLP.n9 VCLP.t26 1363.89
R10742 VCLP.n7 VCLP.t0 1363.89
R10743 VCLP.n5 VCLP.t4 1363.89
R10744 VCLP.n3 VCLP.t22 1363.89
R10745 VCLP.n1 VCLP.t5 1363.89
R10746 VCLP.n109 VCLP.t6 1362.14
R10747 VCLP.n107 VCLP.t41 1362.14
R10748 VCLP.n105 VCLP.t107 1362.14
R10749 VCLP.n103 VCLP.t98 1362.14
R10750 VCLP.n101 VCLP.t35 1362.14
R10751 VCLP.n99 VCLP.t1 1362.14
R10752 VCLP.n97 VCLP.t38 1362.14
R10753 VCLP.n95 VCLP.t2 1362.14
R10754 VCLP.n93 VCLP.t49 1362.14
R10755 VCLP.n91 VCLP.t16 1362.14
R10756 VCLP.n89 VCLP.t80 1362.14
R10757 VCLP.n87 VCLP.t91 1362.14
R10758 VCLP.n85 VCLP.t52 1362.14
R10759 VCLP.n83 VCLP.t48 1362.14
R10760 VCLP.n81 VCLP.t69 1362.14
R10761 VCLP.n79 VCLP.t42 1362.14
R10762 VCLP.n61 VCLP.t95 1362.14
R10763 VCLP.n59 VCLP.t18 1362.14
R10764 VCLP.n57 VCLP.t84 1362.14
R10765 VCLP.n55 VCLP.t76 1362.14
R10766 VCLP.n53 VCLP.t12 1362.14
R10767 VCLP.n51 VCLP.t90 1362.14
R10768 VCLP.n49 VCLP.t15 1362.14
R10769 VCLP.n47 VCLP.t93 1362.14
R10770 VCLP.n45 VCLP.t24 1362.14
R10771 VCLP.n43 VCLP.t105 1362.14
R10772 VCLP.n41 VCLP.t53 1362.14
R10773 VCLP.n39 VCLP.t65 1362.14
R10774 VCLP.n37 VCLP.t30 1362.14
R10775 VCLP.n35 VCLP.t21 1362.14
R10776 VCLP.n33 VCLP.t44 1362.14
R10777 VCLP.n31 VCLP.t19 1362.14
R10778 VCLP.n77 VCLP.t32 1360.68
R10779 VCLP.n75 VCLP.t73 1360.68
R10780 VCLP.n73 VCLP.t20 1360.68
R10781 VCLP.n71 VCLP.t14 1360.68
R10782 VCLP.n69 VCLP.t61 1360.68
R10783 VCLP.n67 VCLP.t25 1360.68
R10784 VCLP.n65 VCLP.t68 1360.68
R10785 VCLP.n63 VCLP.t29 1360.68
R10786 VCLP.n30 VCLP.t37 1360.68
R10787 VCLP.n28 VCLP.t74 1360.68
R10788 VCLP.n26 VCLP.t23 1360.68
R10789 VCLP.n24 VCLP.t17 1360.68
R10790 VCLP.n22 VCLP.t67 1360.68
R10791 VCLP.n20 VCLP.t28 1360.68
R10792 VCLP.n18 VCLP.t71 1360.68
R10793 VCLP.n16 VCLP.t33 1360.68
R10794 VCLP.n14 VCLP.t83 1360.68
R10795 VCLP.n12 VCLP.t47 1360.68
R10796 VCLP.n10 VCLP.t111 1360.68
R10797 VCLP.n8 VCLP.t9 1360.68
R10798 VCLP.n6 VCLP.t86 1360.68
R10799 VCLP.n4 VCLP.t79 1360.68
R10800 VCLP.n2 VCLP.t99 1360.68
R10801 VCLP.n0 VCLP.t75 1360.68
R10802 VCLP.n62 VCLP.n30 23.025
R10803 VCLP.n110 VCLP.n78 15.249
R10804 VCLP.n78 VCLP.n62 8.843
R10805 VCLP VCLP.n110 8.169
R10806 VCLP.n110 VCLP.n109 7.748
R10807 VCLP.n78 VCLP.n77 7.748
R10808 VCLP.n62 VCLP.n61 7.748
R10809 VCLP.n82 VCLP.n81 7.733
R10810 VCLP.n84 VCLP.n83 7.733
R10811 VCLP.n34 VCLP.n33 7.733
R10812 VCLP.n36 VCLP.n35 7.733
R10813 VCLP.n3 VCLP.n2 7.733
R10814 VCLP.n5 VCLP.n4 7.733
R10815 VCLP.n86 VCLP.n85 7.706
R10816 VCLP.n88 VCLP.n87 7.706
R10817 VCLP.n38 VCLP.n37 7.706
R10818 VCLP.n40 VCLP.n39 7.706
R10819 VCLP.n7 VCLP.n6 7.706
R10820 VCLP.n9 VCLP.n8 7.706
R10821 VCLP.n90 VCLP.n89 7.688
R10822 VCLP.n92 VCLP.n91 7.688
R10823 VCLP.n94 VCLP.n93 7.688
R10824 VCLP.n96 VCLP.n95 7.688
R10825 VCLP.n98 VCLP.n97 7.688
R10826 VCLP.n100 VCLP.n99 7.688
R10827 VCLP.n106 VCLP.n105 7.688
R10828 VCLP.n64 VCLP.n63 7.688
R10829 VCLP.n66 VCLP.n65 7.688
R10830 VCLP.n68 VCLP.n67 7.688
R10831 VCLP.n74 VCLP.n73 7.688
R10832 VCLP.n42 VCLP.n41 7.688
R10833 VCLP.n44 VCLP.n43 7.688
R10834 VCLP.n46 VCLP.n45 7.688
R10835 VCLP.n48 VCLP.n47 7.688
R10836 VCLP.n50 VCLP.n49 7.688
R10837 VCLP.n52 VCLP.n51 7.688
R10838 VCLP.n58 VCLP.n57 7.688
R10839 VCLP.n11 VCLP.n10 7.688
R10840 VCLP.n13 VCLP.n12 7.688
R10841 VCLP.n15 VCLP.n14 7.688
R10842 VCLP.n17 VCLP.n16 7.688
R10843 VCLP.n19 VCLP.n18 7.688
R10844 VCLP.n21 VCLP.n20 7.688
R10845 VCLP.n27 VCLP.n26 7.688
R10846 VCLP.n102 VCLP.n101 7.679
R10847 VCLP.n104 VCLP.n103 7.679
R10848 VCLP.n70 VCLP.n69 7.679
R10849 VCLP.n72 VCLP.n71 7.679
R10850 VCLP.n54 VCLP.n53 7.679
R10851 VCLP.n56 VCLP.n55 7.679
R10852 VCLP.n23 VCLP.n22 7.679
R10853 VCLP.n25 VCLP.n24 7.679
R10854 VCLP.n108 VCLP.n107 7.403
R10855 VCLP.n76 VCLP.n75 7.403
R10856 VCLP.n60 VCLP.n59 7.403
R10857 VCLP.n29 VCLP.n28 7.403
R10858 VCLP.n80 VCLP.n79 5.179
R10859 VCLP.n32 VCLP.n31 5.179
R10860 VCLP.n1 VCLP.n0 5.179
R10861 VCLP.n81 VCLP.n80 2.617
R10862 VCLP.n83 VCLP.n82 2.617
R10863 VCLP.n85 VCLP.n84 2.617
R10864 VCLP.n87 VCLP.n86 2.617
R10865 VCLP.n89 VCLP.n88 2.617
R10866 VCLP.n91 VCLP.n90 2.617
R10867 VCLP.n93 VCLP.n92 2.617
R10868 VCLP.n95 VCLP.n94 2.617
R10869 VCLP.n97 VCLP.n96 2.617
R10870 VCLP.n99 VCLP.n98 2.617
R10871 VCLP.n101 VCLP.n100 2.617
R10872 VCLP.n103 VCLP.n102 2.617
R10873 VCLP.n105 VCLP.n104 2.617
R10874 VCLP.n107 VCLP.n106 2.617
R10875 VCLP.n109 VCLP.n108 2.617
R10876 VCLP.n65 VCLP.n64 2.617
R10877 VCLP.n67 VCLP.n66 2.617
R10878 VCLP.n69 VCLP.n68 2.617
R10879 VCLP.n71 VCLP.n70 2.617
R10880 VCLP.n73 VCLP.n72 2.617
R10881 VCLP.n75 VCLP.n74 2.617
R10882 VCLP.n77 VCLP.n76 2.617
R10883 VCLP.n33 VCLP.n32 2.617
R10884 VCLP.n35 VCLP.n34 2.617
R10885 VCLP.n37 VCLP.n36 2.617
R10886 VCLP.n39 VCLP.n38 2.617
R10887 VCLP.n41 VCLP.n40 2.617
R10888 VCLP.n43 VCLP.n42 2.617
R10889 VCLP.n45 VCLP.n44 2.617
R10890 VCLP.n47 VCLP.n46 2.617
R10891 VCLP.n49 VCLP.n48 2.617
R10892 VCLP.n51 VCLP.n50 2.617
R10893 VCLP.n53 VCLP.n52 2.617
R10894 VCLP.n55 VCLP.n54 2.617
R10895 VCLP.n57 VCLP.n56 2.617
R10896 VCLP.n59 VCLP.n58 2.617
R10897 VCLP.n61 VCLP.n60 2.617
R10898 VCLP.n2 VCLP.n1 2.617
R10899 VCLP.n4 VCLP.n3 2.617
R10900 VCLP.n6 VCLP.n5 2.617
R10901 VCLP.n8 VCLP.n7 2.617
R10902 VCLP.n10 VCLP.n9 2.617
R10903 VCLP.n12 VCLP.n11 2.617
R10904 VCLP.n14 VCLP.n13 2.617
R10905 VCLP.n16 VCLP.n15 2.617
R10906 VCLP.n18 VCLP.n17 2.617
R10907 VCLP.n20 VCLP.n19 2.617
R10908 VCLP.n22 VCLP.n21 2.617
R10909 VCLP.n24 VCLP.n23 2.617
R10910 VCLP.n26 VCLP.n25 2.617
R10911 VCLP.n28 VCLP.n27 2.617
R10912 VCLP.n30 VCLP.n29 2.617
R10913 a_9475_n4470.n0 a_9475_n4470.t0 63.08
R10914 a_9475_n4470.n0 a_9475_n4470.t2 41.305
R10915 a_9475_n4470.t1 a_9475_n4470.n0 2.251
R10916 a_9613_n4470.t0 a_9613_n4470.t1 68.741
R10917 a_2049_n7825.t0 a_2049_n7825.t1 42.705
R10918 a_2084_n8026.n0 a_2084_n8026.t0 65.063
R10919 a_2084_n8026.n0 a_2084_n8026.t2 42.011
R10920 a_2084_n8026.t1 a_2084_n8026.n0 2.113
R10921 a_4393_n2422.n3 a_4393_n2422.t2 475.39
R10922 a_4393_n2422.n3 a_4393_n2422.n2 466.481
R10923 a_4393_n2422.t6 a_4393_n2422.t4 228.696
R10924 a_4393_n2422.n2 a_4393_n2422.t1 185.704
R10925 a_4393_n2422.n0 a_4393_n2422.t6 126.761
R10926 a_4393_n2422.n1 a_4393_n2422.t7 126.284
R10927 a_4393_n2422.n1 a_4393_n2422.t0 126.284
R10928 a_4393_n2422.t3 a_4393_n2422.n3 124.375
R10929 a_4393_n2422.t0 a_4393_n2422.n0 115.122
R10930 a_4393_n2422.n0 a_4393_n2422.t5 111.229
R10931 a_4393_n2422.n2 a_4393_n2422.n1 8.764
R10932 a_4413_n7825.t0 a_4413_n7825.t1 42.705
R10933 a_6697_3425.n0 a_6697_3425.t1 358.166
R10934 a_6697_3425.t5 a_6697_3425.t3 337.399
R10935 a_6697_3425.t3 a_6697_3425.t4 285.986
R10936 a_6697_3425.n0 a_6697_3425.t5 282.573
R10937 a_6697_3425.n1 a_6697_3425.t2 202.857
R10938 a_6697_3425.n1 a_6697_3425.n0 173.817
R10939 a_6697_3425.n1 a_6697_3425.t0 20.826
R10940 a_6697_3425.n2 a_6697_3425.n1 20.689
R10941 a_6602_3410.n0 a_6602_3410.t2 362.857
R10942 a_6602_3410.t5 a_6602_3410.t4 337.399
R10943 a_6602_3410.t4 a_6602_3410.t3 298.839
R10944 a_6602_3410.n0 a_6602_3410.t5 280.405
R10945 a_6602_3410.n1 a_6602_3410.t0 200
R10946 a_6602_3410.n1 a_6602_3410.n0 172.311
R10947 a_6602_3410.n2 a_6602_3410.n1 24
R10948 a_6602_3410.n1 a_6602_3410.t1 21.212
R10949 RWL[10].n0 RWL[10].t6 154.243
R10950 RWL[10].n14 RWL[10].t12 149.249
R10951 RWL[10].n13 RWL[10].t1 149.249
R10952 RWL[10].n12 RWL[10].t8 149.249
R10953 RWL[10].n11 RWL[10].t13 149.249
R10954 RWL[10].n10 RWL[10].t10 149.249
R10955 RWL[10].n9 RWL[10].t2 149.249
R10956 RWL[10].n8 RWL[10].t9 149.249
R10957 RWL[10].n7 RWL[10].t15 149.249
R10958 RWL[10].n6 RWL[10].t11 149.249
R10959 RWL[10].n5 RWL[10].t5 149.249
R10960 RWL[10].n4 RWL[10].t14 149.249
R10961 RWL[10].n3 RWL[10].t3 149.249
R10962 RWL[10].n2 RWL[10].t4 149.249
R10963 RWL[10].n1 RWL[10].t7 149.249
R10964 RWL[10].n0 RWL[10].t0 149.249
R10965 RWL[10] RWL[10].n14 42.872
R10966 RWL[10].n1 RWL[10].n0 4.994
R10967 RWL[10].n2 RWL[10].n1 4.994
R10968 RWL[10].n3 RWL[10].n2 4.994
R10969 RWL[10].n4 RWL[10].n3 4.994
R10970 RWL[10].n5 RWL[10].n4 4.994
R10971 RWL[10].n6 RWL[10].n5 4.994
R10972 RWL[10].n7 RWL[10].n6 4.994
R10973 RWL[10].n8 RWL[10].n7 4.994
R10974 RWL[10].n9 RWL[10].n8 4.994
R10975 RWL[10].n10 RWL[10].n9 4.994
R10976 RWL[10].n11 RWL[10].n10 4.994
R10977 RWL[10].n12 RWL[10].n11 4.994
R10978 RWL[10].n13 RWL[10].n12 4.994
R10979 RWL[10].n14 RWL[10].n13 4.994
R10980 a_8340_1216.t0 a_8340_1216.t1 242.857
R10981 a_947_452.n0 a_947_452.t1 358.166
R10982 a_947_452.t5 a_947_452.t4 337.399
R10983 a_947_452.t4 a_947_452.t3 285.986
R10984 a_947_452.n0 a_947_452.t5 282.573
R10985 a_947_452.n1 a_947_452.t0 202.857
R10986 a_947_452.n1 a_947_452.n0 173.817
R10987 a_947_452.n1 a_947_452.t2 20.826
R10988 a_947_452.n2 a_947_452.n1 20.689
R10989 a_1317_452.t0 a_1317_452.t1 242.857
R10990 a_5452_2647.n0 a_5452_2647.t0 362.857
R10991 a_5452_2647.t4 a_5452_2647.t5 337.399
R10992 a_5452_2647.t5 a_5452_2647.t3 298.839
R10993 a_5452_2647.n0 a_5452_2647.t4 280.405
R10994 a_5452_2647.n1 a_5452_2647.t2 200
R10995 a_5452_2647.n1 a_5452_2647.n0 172.311
R10996 a_5452_2647.n2 a_5452_2647.n1 24
R10997 a_5452_2647.n1 a_5452_2647.t1 21.212
R10998 a_5465_2662.t0 a_5465_2662.t1 242.857
R10999 ADC13_OUT[2].n0 ADC13_OUT[2].t4 1354.27
R11000 ADC13_OUT[2].n0 ADC13_OUT[2].t3 821.954
R11001 ADC13_OUT[2].n3 ADC13_OUT[2].t2 327.562
R11002 ADC13_OUT[2].n2 ADC13_OUT[2].t1 266.575
R11003 ADC13_OUT[2].n1 ADC13_OUT[2].n0 149.035
R11004 ADC13_OUT[2].n3 ADC13_OUT[2].n2 56.47
R11005 ADC13_OUT[2].n1 ADC13_OUT[2].t0 46.723
R11006 ADC13_OUT[2] ADC13_OUT[2].n3 38.28
R11007 ADC13_OUT[2].n2 ADC13_OUT[2].n1 17.317
R11008 WWLD[3].n0 WWLD[3].t5 262.032
R11009 WWLD[3].n29 WWLD[3].t8 260.715
R11010 WWLD[3].n27 WWLD[3].t11 260.715
R11011 WWLD[3].n25 WWLD[3].t25 260.715
R11012 WWLD[3].n23 WWLD[3].t19 260.715
R11013 WWLD[3].n21 WWLD[3].t31 260.715
R11014 WWLD[3].n19 WWLD[3].t16 260.715
R11015 WWLD[3].n17 WWLD[3].t7 260.715
R11016 WWLD[3].n15 WWLD[3].t22 260.715
R11017 WWLD[3].n13 WWLD[3].t12 260.715
R11018 WWLD[3].n11 WWLD[3].t20 260.715
R11019 WWLD[3].n9 WWLD[3].t9 260.715
R11020 WWLD[3].n7 WWLD[3].t23 260.715
R11021 WWLD[3].n5 WWLD[3].t17 260.715
R11022 WWLD[3].n3 WWLD[3].t0 260.715
R11023 WWLD[3].n1 WWLD[3].t13 260.715
R11024 WWLD[3].n30 WWLD[3].t24 259.254
R11025 WWLD[3].n28 WWLD[3].t30 259.254
R11026 WWLD[3].n26 WWLD[3].t10 259.254
R11027 WWLD[3].n24 WWLD[3].t26 259.254
R11028 WWLD[3].n22 WWLD[3].t18 259.254
R11029 WWLD[3].n20 WWLD[3].t1 259.254
R11030 WWLD[3].n18 WWLD[3].t14 259.254
R11031 WWLD[3].n16 WWLD[3].t28 259.254
R11032 WWLD[3].n14 WWLD[3].t21 259.254
R11033 WWLD[3].n12 WWLD[3].t4 259.254
R11034 WWLD[3].n10 WWLD[3].t27 259.254
R11035 WWLD[3].n8 WWLD[3].t2 259.254
R11036 WWLD[3].n6 WWLD[3].t3 259.254
R11037 WWLD[3].n4 WWLD[3].t6 259.254
R11038 WWLD[3].n2 WWLD[3].t29 259.254
R11039 WWLD[3].n0 WWLD[3].t15 259.254
R11040 WWLD[3] WWLD[3].n30 44.647
R11041 WWLD[3].n1 WWLD[3].n0 3.576
R11042 WWLD[3].n3 WWLD[3].n2 3.576
R11043 WWLD[3].n5 WWLD[3].n4 3.576
R11044 WWLD[3].n7 WWLD[3].n6 3.576
R11045 WWLD[3].n9 WWLD[3].n8 3.576
R11046 WWLD[3].n11 WWLD[3].n10 3.576
R11047 WWLD[3].n13 WWLD[3].n12 3.576
R11048 WWLD[3].n15 WWLD[3].n14 3.576
R11049 WWLD[3].n17 WWLD[3].n16 3.576
R11050 WWLD[3].n19 WWLD[3].n18 3.576
R11051 WWLD[3].n21 WWLD[3].n20 3.576
R11052 WWLD[3].n23 WWLD[3].n22 3.576
R11053 WWLD[3].n25 WWLD[3].n24 3.576
R11054 WWLD[3].n27 WWLD[3].n26 3.576
R11055 WWLD[3].n29 WWLD[3].n28 3.576
R11056 WWLD[3].n2 WWLD[3].n1 1.317
R11057 WWLD[3].n4 WWLD[3].n3 1.317
R11058 WWLD[3].n6 WWLD[3].n5 1.317
R11059 WWLD[3].n8 WWLD[3].n7 1.317
R11060 WWLD[3].n10 WWLD[3].n9 1.317
R11061 WWLD[3].n12 WWLD[3].n11 1.317
R11062 WWLD[3].n14 WWLD[3].n13 1.317
R11063 WWLD[3].n16 WWLD[3].n15 1.317
R11064 WWLD[3].n18 WWLD[3].n17 1.317
R11065 WWLD[3].n20 WWLD[3].n19 1.317
R11066 WWLD[3].n22 WWLD[3].n21 1.317
R11067 WWLD[3].n24 WWLD[3].n23 1.317
R11068 WWLD[3].n26 WWLD[3].n25 1.317
R11069 WWLD[3].n28 WWLD[3].n27 1.317
R11070 WWLD[3].n30 WWLD[3].n29 1.317
R11071 a_8020_4887.n25 a_8020_4887.t27 561.971
R11072 a_8020_4887.n0 a_8020_4887.t21 449.944
R11073 a_8020_4887.t25 a_8020_4887.n25 108.636
R11074 a_8020_4887.n0 a_8020_4887.t20 74.821
R11075 a_8020_4887.n24 a_8020_4887.t22 63.519
R11076 a_8020_4887.n23 a_8020_4887.t6 63.519
R11077 a_8020_4887.n22 a_8020_4887.t3 63.519
R11078 a_8020_4887.n21 a_8020_4887.t16 63.519
R11079 a_8020_4887.n20 a_8020_4887.t9 63.519
R11080 a_8020_4887.n19 a_8020_4887.t17 63.519
R11081 a_8020_4887.n18 a_8020_4887.t19 63.519
R11082 a_8020_4887.n17 a_8020_4887.t14 63.519
R11083 a_8020_4887.n16 a_8020_4887.t26 63.519
R11084 a_8020_4887.n15 a_8020_4887.t4 63.519
R11085 a_8020_4887.n14 a_8020_4887.t13 63.519
R11086 a_8020_4887.n13 a_8020_4887.t11 63.519
R11087 a_8020_4887.n12 a_8020_4887.t0 63.519
R11088 a_8020_4887.n11 a_8020_4887.t12 63.519
R11089 a_8020_4887.n10 a_8020_4887.t2 63.519
R11090 a_8020_4887.n9 a_8020_4887.t8 63.519
R11091 a_8020_4887.n8 a_8020_4887.t7 63.519
R11092 a_8020_4887.n7 a_8020_4887.t23 63.519
R11093 a_8020_4887.n6 a_8020_4887.t1 63.519
R11094 a_8020_4887.n5 a_8020_4887.t24 63.519
R11095 a_8020_4887.n4 a_8020_4887.t5 63.519
R11096 a_8020_4887.n3 a_8020_4887.t10 63.519
R11097 a_8020_4887.n2 a_8020_4887.t15 63.519
R11098 a_8020_4887.n1 a_8020_4887.t18 63.519
R11099 a_8020_4887.n1 a_8020_4887.n0 8.619
R11100 a_8020_4887.n25 a_8020_4887.n24 2.946
R11101 a_8020_4887.n23 a_8020_4887.n22 2.524
R11102 a_8020_4887.n3 a_8020_4887.n2 2.498
R11103 a_8020_4887.n17 a_8020_4887.n16 2.364
R11104 a_8020_4887.n9 a_8020_4887.n8 2.355
R11105 a_8020_4887.n24 a_8020_4887.n23 1.998
R11106 a_8020_4887.n22 a_8020_4887.n21 1.998
R11107 a_8020_4887.n21 a_8020_4887.n20 1.998
R11108 a_8020_4887.n20 a_8020_4887.n19 1.998
R11109 a_8020_4887.n19 a_8020_4887.n18 1.998
R11110 a_8020_4887.n18 a_8020_4887.n17 1.998
R11111 a_8020_4887.n16 a_8020_4887.n15 1.998
R11112 a_8020_4887.n15 a_8020_4887.n14 1.998
R11113 a_8020_4887.n14 a_8020_4887.n13 1.998
R11114 a_8020_4887.n13 a_8020_4887.n12 1.998
R11115 a_8020_4887.n12 a_8020_4887.n11 1.998
R11116 a_8020_4887.n11 a_8020_4887.n10 1.998
R11117 a_8020_4887.n10 a_8020_4887.n9 1.998
R11118 a_8020_4887.n8 a_8020_4887.n7 1.998
R11119 a_8020_4887.n7 a_8020_4887.n6 1.998
R11120 a_8020_4887.n6 a_8020_4887.n5 1.998
R11121 a_8020_4887.n5 a_8020_4887.n4 1.998
R11122 a_8020_4887.n4 a_8020_4887.n3 1.998
R11123 a_8020_4887.n2 a_8020_4887.n1 1.998
R11124 a_7752_3892.n0 a_7752_3892.t1 362.857
R11125 a_7752_3892.t3 a_7752_3892.t4 337.399
R11126 a_7752_3892.t4 a_7752_3892.t5 298.839
R11127 a_7752_3892.n0 a_7752_3892.t3 280.405
R11128 a_7752_3892.n1 a_7752_3892.t0 200
R11129 a_7752_3892.n1 a_7752_3892.n0 172.311
R11130 a_7752_3892.n2 a_7752_3892.n1 24
R11131 a_7752_3892.n1 a_7752_3892.t2 21.212
R11132 RWL[0].n0 RWL[0].t10 154.243
R11133 RWL[0].n14 RWL[0].t0 149.249
R11134 RWL[0].n13 RWL[0].t5 149.249
R11135 RWL[0].n12 RWL[0].t12 149.249
R11136 RWL[0].n11 RWL[0].t1 149.249
R11137 RWL[0].n10 RWL[0].t14 149.249
R11138 RWL[0].n9 RWL[0].t6 149.249
R11139 RWL[0].n8 RWL[0].t13 149.249
R11140 RWL[0].n7 RWL[0].t3 149.249
R11141 RWL[0].n6 RWL[0].t15 149.249
R11142 RWL[0].n5 RWL[0].t9 149.249
R11143 RWL[0].n4 RWL[0].t2 149.249
R11144 RWL[0].n3 RWL[0].t7 149.249
R11145 RWL[0].n2 RWL[0].t8 149.249
R11146 RWL[0].n1 RWL[0].t11 149.249
R11147 RWL[0].n0 RWL[0].t4 149.249
R11148 RWL[0] RWL[0].n14 42.872
R11149 RWL[0].n1 RWL[0].n0 4.994
R11150 RWL[0].n2 RWL[0].n1 4.994
R11151 RWL[0].n3 RWL[0].n2 4.994
R11152 RWL[0].n4 RWL[0].n3 4.994
R11153 RWL[0].n5 RWL[0].n4 4.994
R11154 RWL[0].n6 RWL[0].n5 4.994
R11155 RWL[0].n7 RWL[0].n6 4.994
R11156 RWL[0].n8 RWL[0].n7 4.994
R11157 RWL[0].n9 RWL[0].n8 4.994
R11158 RWL[0].n10 RWL[0].n9 4.994
R11159 RWL[0].n11 RWL[0].n10 4.994
R11160 RWL[0].n12 RWL[0].n11 4.994
R11161 RWL[0].n13 RWL[0].n12 4.994
R11162 RWL[0].n14 RWL[0].n13 4.994
R11163 a_290_3666.t0 a_290_3666.t1 242.857
R11164 a_290_n953.t35 a_290_n953.n46 171.498
R11165 a_290_n953.n22 a_290_n953.t3 67.378
R11166 a_290_n953.n0 a_290_n953.t16 66.92
R11167 a_290_n953.n1 a_290_n953.t11 66.92
R11168 a_290_n953.n2 a_290_n953.t9 66.92
R11169 a_290_n953.n3 a_290_n953.t18 66.92
R11170 a_290_n953.n4 a_290_n953.t2 66.92
R11171 a_290_n953.n5 a_290_n953.t1 66.92
R11172 a_290_n953.n6 a_290_n953.t40 66.92
R11173 a_290_n953.n7 a_290_n953.t44 66.92
R11174 a_290_n953.n8 a_290_n953.t24 66.92
R11175 a_290_n953.n9 a_290_n953.t29 66.92
R11176 a_290_n953.n10 a_290_n953.t19 66.92
R11177 a_290_n953.n11 a_290_n953.t31 66.92
R11178 a_290_n953.n12 a_290_n953.t23 66.92
R11179 a_290_n953.n13 a_290_n953.t32 66.92
R11180 a_290_n953.n14 a_290_n953.t48 66.92
R11181 a_290_n953.n15 a_290_n953.t46 66.92
R11182 a_290_n953.n16 a_290_n953.t42 66.92
R11183 a_290_n953.n17 a_290_n953.t0 66.92
R11184 a_290_n953.n18 a_290_n953.t22 66.92
R11185 a_290_n953.n19 a_290_n953.t26 66.92
R11186 a_290_n953.n20 a_290_n953.t12 66.92
R11187 a_290_n953.n21 a_290_n953.t15 66.92
R11188 a_290_n953.n22 a_290_n953.t14 66.92
R11189 a_290_n953.n23 a_290_n953.t6 65.518
R11190 a_290_n953.n45 a_290_n953.t5 63.519
R11191 a_290_n953.n44 a_290_n953.t13 63.519
R11192 a_290_n953.n43 a_290_n953.t10 63.519
R11193 a_290_n953.n42 a_290_n953.t4 63.519
R11194 a_290_n953.n41 a_290_n953.t36 63.519
R11195 a_290_n953.n40 a_290_n953.t39 63.519
R11196 a_290_n953.n39 a_290_n953.t21 63.519
R11197 a_290_n953.n38 a_290_n953.t20 63.519
R11198 a_290_n953.n37 a_290_n953.t43 63.519
R11199 a_290_n953.n36 a_290_n953.t38 63.519
R11200 a_290_n953.n35 a_290_n953.t30 63.519
R11201 a_290_n953.n34 a_290_n953.t28 63.519
R11202 a_290_n953.n33 a_290_n953.t33 63.519
R11203 a_290_n953.n32 a_290_n953.t41 63.519
R11204 a_290_n953.n31 a_290_n953.t47 63.519
R11205 a_290_n953.n30 a_290_n953.t37 63.519
R11206 a_290_n953.n29 a_290_n953.t34 63.519
R11207 a_290_n953.n28 a_290_n953.t45 63.519
R11208 a_290_n953.n27 a_290_n953.t27 63.519
R11209 a_290_n953.n26 a_290_n953.t25 63.519
R11210 a_290_n953.n25 a_290_n953.t17 63.519
R11211 a_290_n953.n24 a_290_n953.t7 63.519
R11212 a_290_n953.n23 a_290_n953.t8 63.519
R11213 a_290_n953.n46 a_290_n953.n0 19.59
R11214 a_290_n953.n46 a_290_n953.n45 15.679
R11215 a_290_n953.n44 a_290_n953.n43 2.524
R11216 a_290_n953.n24 a_290_n953.n23 2.498
R11217 a_290_n953.n21 a_290_n953.n22 2.495
R11218 a_290_n953.n1 a_290_n953.n2 2.459
R11219 a_290_n953.n38 a_290_n953.n37 2.364
R11220 a_290_n953.n30 a_290_n953.n29 2.355
R11221 a_290_n953.n7 a_290_n953.n8 2.299
R11222 a_290_n953.n15 a_290_n953.n16 2.29
R11223 a_290_n953.n16 a_290_n953.n17 2.057
R11224 a_290_n953.n8 a_290_n953.n9 2.057
R11225 a_290_n953.n2 a_290_n953.n3 2.057
R11226 a_290_n953.n0 a_290_n953.n1 2.057
R11227 a_290_n953.n45 a_290_n953.n44 1.998
R11228 a_290_n953.n43 a_290_n953.n42 1.998
R11229 a_290_n953.n42 a_290_n953.n41 1.998
R11230 a_290_n953.n41 a_290_n953.n40 1.998
R11231 a_290_n953.n40 a_290_n953.n39 1.998
R11232 a_290_n953.n39 a_290_n953.n38 1.998
R11233 a_290_n953.n37 a_290_n953.n36 1.998
R11234 a_290_n953.n36 a_290_n953.n35 1.998
R11235 a_290_n953.n35 a_290_n953.n34 1.998
R11236 a_290_n953.n34 a_290_n953.n33 1.998
R11237 a_290_n953.n33 a_290_n953.n32 1.998
R11238 a_290_n953.n32 a_290_n953.n31 1.998
R11239 a_290_n953.n31 a_290_n953.n30 1.998
R11240 a_290_n953.n29 a_290_n953.n28 1.998
R11241 a_290_n953.n28 a_290_n953.n27 1.998
R11242 a_290_n953.n27 a_290_n953.n26 1.998
R11243 a_290_n953.n26 a_290_n953.n25 1.998
R11244 a_290_n953.n25 a_290_n953.n24 1.998
R11245 a_290_n953.n20 a_290_n953.n21 1.995
R11246 a_290_n953.n19 a_290_n953.n20 1.995
R11247 a_290_n953.n18 a_290_n953.n19 1.995
R11248 a_290_n953.n17 a_290_n953.n18 1.995
R11249 a_290_n953.n14 a_290_n953.n15 1.995
R11250 a_290_n953.n13 a_290_n953.n14 1.995
R11251 a_290_n953.n12 a_290_n953.n13 1.995
R11252 a_290_n953.n11 a_290_n953.n12 1.995
R11253 a_290_n953.n10 a_290_n953.n11 1.995
R11254 a_290_n953.n9 a_290_n953.n10 1.995
R11255 a_290_n953.n6 a_290_n953.n7 1.995
R11256 a_290_n953.n5 a_290_n953.n6 1.995
R11257 a_290_n953.n4 a_290_n953.n5 1.995
R11258 a_290_n953.n3 a_290_n953.n4 1.995
R11259 a_6602_2165.n0 a_6602_2165.t1 362.857
R11260 a_6602_2165.t3 a_6602_2165.t5 337.399
R11261 a_6602_2165.t5 a_6602_2165.t4 298.839
R11262 a_6602_2165.n0 a_6602_2165.t3 280.405
R11263 a_6602_2165.n1 a_6602_2165.t2 200
R11264 a_6602_2165.n1 a_6602_2165.n0 172.311
R11265 a_6602_2165.n2 a_6602_2165.n1 24
R11266 a_6602_2165.n1 a_6602_2165.t0 21.212
R11267 a_6697_2180.n0 a_6697_2180.t1 358.166
R11268 a_6697_2180.t5 a_6697_2180.t3 337.399
R11269 a_6697_2180.t3 a_6697_2180.t4 285.986
R11270 a_6697_2180.n0 a_6697_2180.t5 282.573
R11271 a_6697_2180.n1 a_6697_2180.t2 202.857
R11272 a_6697_2180.n1 a_6697_2180.n0 173.817
R11273 a_6697_2180.n1 a_6697_2180.t0 20.826
R11274 a_6697_2180.n2 a_6697_2180.n1 20.689
R11275 a_865_1216.t0 a_865_1216.t1 242.857
R11276 a_947_4445.n0 a_947_4445.t2 358.166
R11277 a_947_4445.t5 a_947_4445.t3 337.399
R11278 a_947_4445.t3 a_947_4445.t4 285.986
R11279 a_947_4445.n0 a_947_4445.t5 282.573
R11280 a_947_4445.n1 a_947_4445.t1 202.857
R11281 a_947_4445.n1 a_947_4445.n0 173.817
R11282 a_947_4445.n1 a_947_4445.t0 20.826
R11283 a_947_4445.n2 a_947_4445.n1 20.689
R11284 a_852_4430.n0 a_852_4430.t1 362.857
R11285 a_852_4430.t3 a_852_4430.t4 337.399
R11286 a_852_4430.t4 a_852_4430.t5 298.839
R11287 a_852_4430.n0 a_852_4430.t3 280.405
R11288 a_852_4430.n1 a_852_4430.t2 200
R11289 a_852_4430.n1 a_852_4430.n0 172.311
R11290 a_852_4430.n2 a_852_4430.n1 24
R11291 a_852_4430.n1 a_852_4430.t0 21.212
R11292 a_3822_3666.n0 a_3822_3666.t0 358.166
R11293 a_3822_3666.t5 a_3822_3666.t4 337.399
R11294 a_3822_3666.t4 a_3822_3666.t3 285.986
R11295 a_3822_3666.n0 a_3822_3666.t5 282.573
R11296 a_3822_3666.n1 a_3822_3666.t2 202.857
R11297 a_3822_3666.n1 a_3822_3666.n0 173.817
R11298 a_3822_3666.n1 a_3822_3666.t1 20.826
R11299 a_3822_3666.n2 a_3822_3666.n1 20.689
R11300 a_4192_3666.t0 a_4192_3666.t1 242.857
R11301 a_4397_1216.n0 a_4397_1216.t1 358.166
R11302 a_4397_1216.t4 a_4397_1216.t5 337.399
R11303 a_4397_1216.t5 a_4397_1216.t3 285.986
R11304 a_4397_1216.n0 a_4397_1216.t4 282.573
R11305 a_4397_1216.n1 a_4397_1216.t2 202.857
R11306 a_4397_1216.n1 a_4397_1216.n0 173.817
R11307 a_4397_1216.n1 a_4397_1216.t0 20.826
R11308 a_4397_1216.n2 a_4397_1216.n1 20.689
R11309 a_4767_1216.t0 a_4767_1216.t1 242.857
R11310 WWL[7].n0 WWL[7].t25 262.032
R11311 WWL[7].n29 WWL[7].t28 260.715
R11312 WWL[7].n27 WWL[7].t31 260.715
R11313 WWL[7].n25 WWL[7].t12 260.715
R11314 WWL[7].n23 WWL[7].t7 260.715
R11315 WWL[7].n21 WWL[7].t17 260.715
R11316 WWL[7].n19 WWL[7].t3 260.715
R11317 WWL[7].n17 WWL[7].t27 260.715
R11318 WWL[7].n15 WWL[7].t10 260.715
R11319 WWL[7].n13 WWL[7].t0 260.715
R11320 WWL[7].n11 WWL[7].t8 260.715
R11321 WWL[7].n9 WWL[7].t29 260.715
R11322 WWL[7].n7 WWL[7].t11 260.715
R11323 WWL[7].n5 WWL[7].t5 260.715
R11324 WWL[7].n3 WWL[7].t20 260.715
R11325 WWL[7].n1 WWL[7].t1 260.715
R11326 WWL[7].n30 WWL[7].t13 259.254
R11327 WWL[7].n28 WWL[7].t19 259.254
R11328 WWL[7].n26 WWL[7].t30 259.254
R11329 WWL[7].n24 WWL[7].t14 259.254
R11330 WWL[7].n22 WWL[7].t6 259.254
R11331 WWL[7].n20 WWL[7].t21 259.254
R11332 WWL[7].n18 WWL[7].t2 259.254
R11333 WWL[7].n16 WWL[7].t16 259.254
R11334 WWL[7].n14 WWL[7].t9 259.254
R11335 WWL[7].n12 WWL[7].t24 259.254
R11336 WWL[7].n10 WWL[7].t15 259.254
R11337 WWL[7].n8 WWL[7].t22 259.254
R11338 WWL[7].n6 WWL[7].t23 259.254
R11339 WWL[7].n4 WWL[7].t26 259.254
R11340 WWL[7].n2 WWL[7].t18 259.254
R11341 WWL[7].n0 WWL[7].t4 259.254
R11342 WWL[7] WWL[7].n30 44.647
R11343 WWL[7].n1 WWL[7].n0 3.576
R11344 WWL[7].n3 WWL[7].n2 3.576
R11345 WWL[7].n5 WWL[7].n4 3.576
R11346 WWL[7].n7 WWL[7].n6 3.576
R11347 WWL[7].n9 WWL[7].n8 3.576
R11348 WWL[7].n11 WWL[7].n10 3.576
R11349 WWL[7].n13 WWL[7].n12 3.576
R11350 WWL[7].n15 WWL[7].n14 3.576
R11351 WWL[7].n17 WWL[7].n16 3.576
R11352 WWL[7].n19 WWL[7].n18 3.576
R11353 WWL[7].n21 WWL[7].n20 3.576
R11354 WWL[7].n23 WWL[7].n22 3.576
R11355 WWL[7].n25 WWL[7].n24 3.576
R11356 WWL[7].n27 WWL[7].n26 3.576
R11357 WWL[7].n29 WWL[7].n28 3.576
R11358 WWL[7].n2 WWL[7].n1 1.317
R11359 WWL[7].n4 WWL[7].n3 1.317
R11360 WWL[7].n6 WWL[7].n5 1.317
R11361 WWL[7].n8 WWL[7].n7 1.317
R11362 WWL[7].n10 WWL[7].n9 1.317
R11363 WWL[7].n12 WWL[7].n11 1.317
R11364 WWL[7].n14 WWL[7].n13 1.317
R11365 WWL[7].n16 WWL[7].n15 1.317
R11366 WWL[7].n18 WWL[7].n17 1.317
R11367 WWL[7].n20 WWL[7].n19 1.317
R11368 WWL[7].n22 WWL[7].n21 1.317
R11369 WWL[7].n24 WWL[7].n23 1.317
R11370 WWL[7].n26 WWL[7].n25 1.317
R11371 WWL[7].n28 WWL[7].n27 1.317
R11372 WWL[7].n30 WWL[7].n29 1.317
R11373 a_5145_4887.n25 a_5145_4887.t27 561.971
R11374 a_5145_4887.n0 a_5145_4887.t20 449.944
R11375 a_5145_4887.t24 a_5145_4887.n25 108.636
R11376 a_5145_4887.n0 a_5145_4887.t19 74.821
R11377 a_5145_4887.n24 a_5145_4887.t25 63.519
R11378 a_5145_4887.n23 a_5145_4887.t6 63.519
R11379 a_5145_4887.n22 a_5145_4887.t2 63.519
R11380 a_5145_4887.n21 a_5145_4887.t16 63.519
R11381 a_5145_4887.n20 a_5145_4887.t9 63.519
R11382 a_5145_4887.n19 a_5145_4887.t17 63.519
R11383 a_5145_4887.n18 a_5145_4887.t21 63.519
R11384 a_5145_4887.n17 a_5145_4887.t14 63.519
R11385 a_5145_4887.n16 a_5145_4887.t26 63.519
R11386 a_5145_4887.n15 a_5145_4887.t3 63.519
R11387 a_5145_4887.n14 a_5145_4887.t13 63.519
R11388 a_5145_4887.n13 a_5145_4887.t10 63.519
R11389 a_5145_4887.n12 a_5145_4887.t5 63.519
R11390 a_5145_4887.n11 a_5145_4887.t12 63.519
R11391 a_5145_4887.n10 a_5145_4887.t1 63.519
R11392 a_5145_4887.n9 a_5145_4887.t8 63.519
R11393 a_5145_4887.n8 a_5145_4887.t7 63.519
R11394 a_5145_4887.n7 a_5145_4887.t22 63.519
R11395 a_5145_4887.n6 a_5145_4887.t0 63.519
R11396 a_5145_4887.n5 a_5145_4887.t23 63.519
R11397 a_5145_4887.n4 a_5145_4887.t4 63.519
R11398 a_5145_4887.n3 a_5145_4887.t11 63.519
R11399 a_5145_4887.n2 a_5145_4887.t15 63.519
R11400 a_5145_4887.n1 a_5145_4887.t18 63.519
R11401 a_5145_4887.n1 a_5145_4887.n0 8.619
R11402 a_5145_4887.n25 a_5145_4887.n24 2.946
R11403 a_5145_4887.n23 a_5145_4887.n22 2.524
R11404 a_5145_4887.n3 a_5145_4887.n2 2.498
R11405 a_5145_4887.n17 a_5145_4887.n16 2.364
R11406 a_5145_4887.n9 a_5145_4887.n8 2.355
R11407 a_5145_4887.n24 a_5145_4887.n23 1.998
R11408 a_5145_4887.n22 a_5145_4887.n21 1.998
R11409 a_5145_4887.n21 a_5145_4887.n20 1.998
R11410 a_5145_4887.n20 a_5145_4887.n19 1.998
R11411 a_5145_4887.n19 a_5145_4887.n18 1.998
R11412 a_5145_4887.n18 a_5145_4887.n17 1.998
R11413 a_5145_4887.n16 a_5145_4887.n15 1.998
R11414 a_5145_4887.n15 a_5145_4887.n14 1.998
R11415 a_5145_4887.n14 a_5145_4887.n13 1.998
R11416 a_5145_4887.n13 a_5145_4887.n12 1.998
R11417 a_5145_4887.n12 a_5145_4887.n11 1.998
R11418 a_5145_4887.n11 a_5145_4887.n10 1.998
R11419 a_5145_4887.n10 a_5145_4887.n9 1.998
R11420 a_5145_4887.n8 a_5145_4887.n7 1.998
R11421 a_5145_4887.n7 a_5145_4887.n6 1.998
R11422 a_5145_4887.n6 a_5145_4887.n5 1.998
R11423 a_5145_4887.n5 a_5145_4887.n4 1.998
R11424 a_5145_4887.n4 a_5145_4887.n3 1.998
R11425 a_5145_4887.n2 a_5145_4887.n1 1.998
R11426 a_4877_1924.n0 a_4877_1924.t2 362.857
R11427 a_4877_1924.t4 a_4877_1924.t3 337.399
R11428 a_4877_1924.t3 a_4877_1924.t5 298.839
R11429 a_4877_1924.n0 a_4877_1924.t4 280.405
R11430 a_4877_1924.n1 a_4877_1924.t0 200
R11431 a_4877_1924.n1 a_4877_1924.n0 172.311
R11432 a_4877_1924.n2 a_4877_1924.n1 24
R11433 a_4877_1924.n1 a_4877_1924.t1 21.212
R11434 a_1427_n527.n0 a_1427_n527.t1 362.857
R11435 a_1427_n527.t4 a_1427_n527.t5 337.399
R11436 a_1427_n527.t5 a_1427_n527.t3 298.839
R11437 a_1427_n527.n0 a_1427_n527.t4 280.405
R11438 a_1427_n527.n1 a_1427_n527.t0 200
R11439 a_1427_n527.n1 a_1427_n527.n0 172.311
R11440 a_1427_n527.n2 a_1427_n527.n1 24
R11441 a_1427_n527.n1 a_1427_n527.t2 21.212
R11442 a_1440_n512.t0 a_1440_n512.t1 242.857
R11443 ADC15_OUT[1].n0 ADC15_OUT[1].t4 1355.37
R11444 ADC15_OUT[1].n0 ADC15_OUT[1].t3 820.859
R11445 ADC15_OUT[1].n3 ADC15_OUT[1].t0 336.667
R11446 ADC15_OUT[1].n2 ADC15_OUT[1].t2 266.644
R11447 ADC15_OUT[1].n1 ADC15_OUT[1].n0 149.035
R11448 ADC15_OUT[1].n3 ADC15_OUT[1].n2 47.435
R11449 ADC15_OUT[1].n1 ADC15_OUT[1].t1 45.968
R11450 ADC15_OUT[1] ADC15_OUT[1].n3 45.82
R11451 ADC15_OUT[1].n2 ADC15_OUT[1].n1 17.317
R11452 a_13864_n5850.n0 a_13864_n5850.t4 1465.51
R11453 a_13864_n5850.n0 a_13864_n5850.t3 712.44
R11454 a_13864_n5850.n1 a_13864_n5850.t0 375.067
R11455 a_13864_n5850.n1 a_13864_n5850.t2 272.668
R11456 a_13864_n5850.n2 a_13864_n5850.n0 143.764
R11457 a_13864_n5850.t1 a_13864_n5850.n2 78.193
R11458 a_13864_n5850.n2 a_13864_n5850.n1 4.517
R11459 SA_OUT[7].n0 SA_OUT[7].t4 661.027
R11460 SA_OUT[7].n0 SA_OUT[7].t3 392.255
R11461 SA_OUT[7].n1 SA_OUT[7].t1 223.716
R11462 SA_OUT[7].n2 SA_OUT[7].t0 153.977
R11463 SA_OUT[7].n1 SA_OUT[7].n0 143.764
R11464 SA_OUT[7].n3 SA_OUT[7].t2 58.354
R11465 SA_OUT[7] SA_OUT[7].n3 15.469
R11466 SA_OUT[7].n2 SA_OUT[7].n1 4.517
R11467 SA_OUT[7].n3 SA_OUT[7].n2 1.505
R11468 a_3822_n512.n0 a_3822_n512.t2 358.166
R11469 a_3822_n512.t4 a_3822_n512.t3 337.399
R11470 a_3822_n512.t3 a_3822_n512.t5 285.986
R11471 a_3822_n512.n0 a_3822_n512.t4 282.573
R11472 a_3822_n512.n1 a_3822_n512.t1 202.857
R11473 a_3822_n512.n1 a_3822_n512.n0 173.817
R11474 a_3822_n512.n1 a_3822_n512.t0 20.826
R11475 a_3822_n512.n2 a_3822_n512.n1 20.689
R11476 a_3727_n527.n0 a_3727_n527.t2 362.857
R11477 a_3727_n527.t4 a_3727_n527.t5 337.399
R11478 a_3727_n527.t5 a_3727_n527.t3 298.839
R11479 a_3727_n527.n0 a_3727_n527.t4 280.405
R11480 a_3727_n527.n1 a_3727_n527.t0 200
R11481 a_3727_n527.n1 a_3727_n527.n0 172.311
R11482 a_3727_n527.n2 a_3727_n527.n1 24
R11483 a_3727_n527.n1 a_3727_n527.t1 21.212
R11484 a_10659_n7203.n0 a_10659_n7203.t0 63.08
R11485 a_10659_n7203.t1 a_10659_n7203.n0 41.306
R11486 a_10659_n7203.n0 a_10659_n7203.t2 2.251
R11487 a_10797_n7203.t1 a_10797_n7203.t0 68.741
R11488 a_8977_n2234.n2 a_8977_n2234.t0 282.97
R11489 a_8977_n2234.n1 a_8977_n2234.t3 240.683
R11490 a_8977_n2234.n0 a_8977_n2234.t4 209.208
R11491 a_8977_n2234.n0 a_8977_n2234.t2 194.167
R11492 a_8977_n2234.t1 a_8977_n2234.n2 183.404
R11493 a_8977_n2234.n1 a_8977_n2234.n0 14.805
R11494 a_8977_n2234.n2 a_8977_n2234.n1 6.415
R11495 a_9100_n2132.n0 a_9100_n2132.t2 489.336
R11496 a_9100_n2132.n0 a_9100_n2132.t1 243.258
R11497 a_9100_n2132.t0 a_9100_n2132.n0 214.415
R11498 a_4972_1216.n0 a_4972_1216.t2 358.166
R11499 a_4972_1216.t4 a_4972_1216.t3 337.399
R11500 a_4972_1216.t3 a_4972_1216.t5 285.986
R11501 a_4972_1216.n0 a_4972_1216.t4 282.573
R11502 a_4972_1216.n1 a_4972_1216.t0 202.857
R11503 a_4972_1216.n1 a_4972_1216.n0 173.817
R11504 a_4972_1216.n1 a_4972_1216.t1 20.826
R11505 a_4972_1216.n2 a_4972_1216.n1 20.689
R11506 a_4877_1201.n0 a_4877_1201.t2 362.857
R11507 a_4877_1201.t4 a_4877_1201.t3 337.399
R11508 a_4877_1201.t3 a_4877_1201.t5 298.839
R11509 a_4877_1201.n0 a_4877_1201.t4 280.405
R11510 a_4877_1201.n1 a_4877_1201.t0 200
R11511 a_4877_1201.n1 a_4877_1201.n0 172.311
R11512 a_4877_1201.n2 a_4877_1201.n1 24
R11513 a_4877_1201.n1 a_4877_1201.t1 21.212
R11514 a_3185_n1371.n1 a_3185_n1371.t3 550.94
R11515 a_3185_n1371.n1 a_3185_n1371.t4 500.621
R11516 a_3185_n1371.t1 a_3185_n1371.n2 192.787
R11517 a_3185_n1371.n0 a_3185_n1371.t0 163.997
R11518 a_3185_n1371.n2 a_3185_n1371.n1 149.035
R11519 a_3185_n1371.n0 a_3185_n1371.t2 54.068
R11520 a_3185_n1371.n2 a_3185_n1371.n0 17.317
R11521 a_7847_3907.n0 a_7847_3907.t2 358.166
R11522 a_7847_3907.t4 a_7847_3907.t5 337.399
R11523 a_7847_3907.t5 a_7847_3907.t3 285.986
R11524 a_7847_3907.n0 a_7847_3907.t4 282.573
R11525 a_7847_3907.n1 a_7847_3907.t0 202.857
R11526 a_7847_3907.n1 a_7847_3907.n0 173.817
R11527 a_7847_3907.n1 a_7847_3907.t1 20.826
R11528 a_7847_3907.n2 a_7847_3907.n1 20.689
R11529 a_8217_3907.t0 a_8217_3907.t1 242.857
R11530 a_3822_975.n0 a_3822_975.t1 358.166
R11531 a_3822_975.t3 a_3822_975.t5 337.399
R11532 a_3822_975.t5 a_3822_975.t4 285.986
R11533 a_3822_975.n0 a_3822_975.t3 282.573
R11534 a_3822_975.n1 a_3822_975.t2 202.857
R11535 a_3822_975.n1 a_3822_975.n0 173.817
R11536 a_3822_975.n1 a_3822_975.t0 20.826
R11537 a_3822_975.n2 a_3822_975.n1 20.689
R11538 a_3727_960.n0 a_3727_960.t1 362.857
R11539 a_3727_960.t4 a_3727_960.t3 337.399
R11540 a_3727_960.t3 a_3727_960.t5 298.839
R11541 a_3727_960.n0 a_3727_960.t4 280.405
R11542 a_3727_960.n1 a_3727_960.t2 200
R11543 a_3727_960.n1 a_3727_960.n0 172.311
R11544 a_3727_960.n2 a_3727_960.n1 24
R11545 a_3727_960.n1 a_3727_960.t0 21.212
R11546 a_4972_n1053.n0 a_4972_n1053.t1 358.166
R11547 a_4972_n1053.t3 a_4972_n1053.t5 337.399
R11548 a_4972_n1053.t5 a_4972_n1053.t4 285.986
R11549 a_4972_n1053.n0 a_4972_n1053.t3 282.573
R11550 a_4972_n1053.n1 a_4972_n1053.t2 202.857
R11551 a_4972_n1053.n1 a_4972_n1053.n0 173.817
R11552 a_4972_n1053.n1 a_4972_n1053.t0 20.826
R11553 a_4972_n1053.n2 a_4972_n1053.n1 20.689
R11554 a_4877_n1068.n0 a_4877_n1068.t1 362.857
R11555 a_4877_n1068.t3 a_4877_n1068.t4 337.399
R11556 a_4877_n1068.t4 a_4877_n1068.t5 298.839
R11557 a_4877_n1068.n0 a_4877_n1068.t3 280.405
R11558 a_4877_n1068.n1 a_4877_n1068.t2 200
R11559 a_4877_n1068.n1 a_4877_n1068.n0 172.311
R11560 a_4877_n1068.n2 a_4877_n1068.n1 24
R11561 a_4877_n1068.n1 a_4877_n1068.t0 21.212
R11562 RWL[2].n0 RWL[2].t9 154.243
R11563 RWL[2].n14 RWL[2].t15 149.249
R11564 RWL[2].n13 RWL[2].t4 149.249
R11565 RWL[2].n12 RWL[2].t11 149.249
R11566 RWL[2].n11 RWL[2].t0 149.249
R11567 RWL[2].n10 RWL[2].t13 149.249
R11568 RWL[2].n9 RWL[2].t5 149.249
R11569 RWL[2].n8 RWL[2].t12 149.249
R11570 RWL[2].n7 RWL[2].t2 149.249
R11571 RWL[2].n6 RWL[2].t14 149.249
R11572 RWL[2].n5 RWL[2].t8 149.249
R11573 RWL[2].n4 RWL[2].t1 149.249
R11574 RWL[2].n3 RWL[2].t6 149.249
R11575 RWL[2].n2 RWL[2].t7 149.249
R11576 RWL[2].n1 RWL[2].t10 149.249
R11577 RWL[2].n0 RWL[2].t3 149.249
R11578 RWL[2] RWL[2].n14 42.872
R11579 RWL[2].n1 RWL[2].n0 4.994
R11580 RWL[2].n2 RWL[2].n1 4.994
R11581 RWL[2].n3 RWL[2].n2 4.994
R11582 RWL[2].n4 RWL[2].n3 4.994
R11583 RWL[2].n5 RWL[2].n4 4.994
R11584 RWL[2].n6 RWL[2].n5 4.994
R11585 RWL[2].n7 RWL[2].n6 4.994
R11586 RWL[2].n8 RWL[2].n7 4.994
R11587 RWL[2].n9 RWL[2].n8 4.994
R11588 RWL[2].n10 RWL[2].n9 4.994
R11589 RWL[2].n11 RWL[2].n10 4.994
R11590 RWL[2].n12 RWL[2].n11 4.994
R11591 RWL[2].n13 RWL[2].n12 4.994
R11592 RWL[2].n14 RWL[2].n13 4.994
R11593 a_2015_3184.t0 a_2015_3184.t1 242.857
R11594 a_2015_n953.t33 a_2015_n953.n46 176.385
R11595 a_2015_n953.n22 a_2015_n953.t13 67.378
R11596 a_2015_n953.n0 a_2015_n953.t15 66.92
R11597 a_2015_n953.n1 a_2015_n953.t6 66.92
R11598 a_2015_n953.n2 a_2015_n953.t11 66.92
R11599 a_2015_n953.n3 a_2015_n953.t9 66.92
R11600 a_2015_n953.n4 a_2015_n953.t0 66.92
R11601 a_2015_n953.n5 a_2015_n953.t48 66.92
R11602 a_2015_n953.n6 a_2015_n953.t39 66.92
R11603 a_2015_n953.n7 a_2015_n953.t42 66.92
R11604 a_2015_n953.n8 a_2015_n953.t21 66.92
R11605 a_2015_n953.n9 a_2015_n953.t27 66.92
R11606 a_2015_n953.n10 a_2015_n953.t17 66.92
R11607 a_2015_n953.n11 a_2015_n953.t29 66.92
R11608 a_2015_n953.n12 a_2015_n953.t25 66.92
R11609 a_2015_n953.n13 a_2015_n953.t30 66.92
R11610 a_2015_n953.n14 a_2015_n953.t47 66.92
R11611 a_2015_n953.n15 a_2015_n953.t45 66.92
R11612 a_2015_n953.n16 a_2015_n953.t46 66.92
R11613 a_2015_n953.n17 a_2015_n953.t23 66.92
R11614 a_2015_n953.n18 a_2015_n953.t20 66.92
R11615 a_2015_n953.n19 a_2015_n953.t24 66.92
R11616 a_2015_n953.n20 a_2015_n953.t7 66.92
R11617 a_2015_n953.n21 a_2015_n953.t3 66.92
R11618 a_2015_n953.n22 a_2015_n953.t12 66.92
R11619 a_2015_n953.n23 a_2015_n953.t1 65.518
R11620 a_2015_n953.n45 a_2015_n953.t2 63.519
R11621 a_2015_n953.n44 a_2015_n953.t10 63.519
R11622 a_2015_n953.n43 a_2015_n953.t14 63.519
R11623 a_2015_n953.n42 a_2015_n953.t16 63.519
R11624 a_2015_n953.n41 a_2015_n953.t34 63.519
R11625 a_2015_n953.n40 a_2015_n953.t38 63.519
R11626 a_2015_n953.n39 a_2015_n953.t19 63.519
R11627 a_2015_n953.n38 a_2015_n953.t18 63.519
R11628 a_2015_n953.n37 a_2015_n953.t41 63.519
R11629 a_2015_n953.n36 a_2015_n953.t37 63.519
R11630 a_2015_n953.n35 a_2015_n953.t28 63.519
R11631 a_2015_n953.n34 a_2015_n953.t31 63.519
R11632 a_2015_n953.n33 a_2015_n953.t35 63.519
R11633 a_2015_n953.n32 a_2015_n953.t40 63.519
R11634 a_2015_n953.n31 a_2015_n953.t43 63.519
R11635 a_2015_n953.n30 a_2015_n953.t36 63.519
R11636 a_2015_n953.n29 a_2015_n953.t32 63.519
R11637 a_2015_n953.n28 a_2015_n953.t44 63.519
R11638 a_2015_n953.n27 a_2015_n953.t26 63.519
R11639 a_2015_n953.n26 a_2015_n953.t22 63.519
R11640 a_2015_n953.n25 a_2015_n953.t8 63.519
R11641 a_2015_n953.n24 a_2015_n953.t4 63.519
R11642 a_2015_n953.n23 a_2015_n953.t5 63.519
R11643 a_2015_n953.n46 a_2015_n953.n45 18.144
R11644 a_2015_n953.n46 a_2015_n953.n0 17.125
R11645 a_2015_n953.n44 a_2015_n953.n43 2.524
R11646 a_2015_n953.n24 a_2015_n953.n23 2.498
R11647 a_2015_n953.n21 a_2015_n953.n22 2.495
R11648 a_2015_n953.n1 a_2015_n953.n2 2.459
R11649 a_2015_n953.n38 a_2015_n953.n37 2.364
R11650 a_2015_n953.n30 a_2015_n953.n29 2.355
R11651 a_2015_n953.n7 a_2015_n953.n8 2.299
R11652 a_2015_n953.n15 a_2015_n953.n16 2.29
R11653 a_2015_n953.n16 a_2015_n953.n17 2.057
R11654 a_2015_n953.n8 a_2015_n953.n9 2.057
R11655 a_2015_n953.n2 a_2015_n953.n3 2.057
R11656 a_2015_n953.n0 a_2015_n953.n1 2.057
R11657 a_2015_n953.n45 a_2015_n953.n44 1.998
R11658 a_2015_n953.n43 a_2015_n953.n42 1.998
R11659 a_2015_n953.n42 a_2015_n953.n41 1.998
R11660 a_2015_n953.n41 a_2015_n953.n40 1.998
R11661 a_2015_n953.n40 a_2015_n953.n39 1.998
R11662 a_2015_n953.n39 a_2015_n953.n38 1.998
R11663 a_2015_n953.n37 a_2015_n953.n36 1.998
R11664 a_2015_n953.n36 a_2015_n953.n35 1.998
R11665 a_2015_n953.n35 a_2015_n953.n34 1.998
R11666 a_2015_n953.n34 a_2015_n953.n33 1.998
R11667 a_2015_n953.n33 a_2015_n953.n32 1.998
R11668 a_2015_n953.n32 a_2015_n953.n31 1.998
R11669 a_2015_n953.n31 a_2015_n953.n30 1.998
R11670 a_2015_n953.n29 a_2015_n953.n28 1.998
R11671 a_2015_n953.n28 a_2015_n953.n27 1.998
R11672 a_2015_n953.n27 a_2015_n953.n26 1.998
R11673 a_2015_n953.n26 a_2015_n953.n25 1.998
R11674 a_2015_n953.n25 a_2015_n953.n24 1.998
R11675 a_2015_n953.n20 a_2015_n953.n21 1.995
R11676 a_2015_n953.n19 a_2015_n953.n20 1.995
R11677 a_2015_n953.n18 a_2015_n953.n19 1.995
R11678 a_2015_n953.n17 a_2015_n953.n18 1.995
R11679 a_2015_n953.n14 a_2015_n953.n15 1.995
R11680 a_2015_n953.n13 a_2015_n953.n14 1.995
R11681 a_2015_n953.n12 a_2015_n953.n13 1.995
R11682 a_2015_n953.n11 a_2015_n953.n12 1.995
R11683 a_2015_n953.n10 a_2015_n953.n11 1.995
R11684 a_2015_n953.n9 a_2015_n953.n10 1.995
R11685 a_2015_n953.n6 a_2015_n953.n7 1.995
R11686 a_2015_n953.n5 a_2015_n953.n6 1.995
R11687 a_2015_n953.n4 a_2015_n953.n5 1.995
R11688 a_2015_n953.n3 a_2015_n953.n4 1.995
R11689 a_2590_n30.t0 a_2590_n30.t1 242.857
R11690 a_4877_2406.n0 a_4877_2406.t2 362.857
R11691 a_4877_2406.t5 a_4877_2406.t4 337.399
R11692 a_4877_2406.t4 a_4877_2406.t3 298.839
R11693 a_4877_2406.n0 a_4877_2406.t5 280.405
R11694 a_4877_2406.n1 a_4877_2406.t0 200
R11695 a_4877_2406.n1 a_4877_2406.n0 172.311
R11696 a_4877_2406.n2 a_4877_2406.n1 24
R11697 a_4877_2406.n1 a_4877_2406.t1 21.212
R11698 a_4890_2421.t0 a_4890_2421.t1 242.857
R11699 a_7177_2406.n0 a_7177_2406.t1 362.857
R11700 a_7177_2406.t3 a_7177_2406.t4 337.399
R11701 a_7177_2406.t4 a_7177_2406.t5 298.839
R11702 a_7177_2406.n0 a_7177_2406.t3 280.405
R11703 a_7177_2406.n1 a_7177_2406.t0 200
R11704 a_7177_2406.n1 a_7177_2406.n0 172.311
R11705 a_7177_2406.n2 a_7177_2406.n1 24
R11706 a_7177_2406.n1 a_7177_2406.t2 21.212
R11707 a_7272_2421.n0 a_7272_2421.t2 358.166
R11708 a_7272_2421.t4 a_7272_2421.t3 337.399
R11709 a_7272_2421.t3 a_7272_2421.t5 285.986
R11710 a_7272_2421.n0 a_7272_2421.t4 282.573
R11711 a_7272_2421.n1 a_7272_2421.t0 202.857
R11712 a_7272_2421.n1 a_7272_2421.n0 173.817
R11713 a_7272_2421.n1 a_7272_2421.t1 20.826
R11714 a_7272_2421.n2 a_7272_2421.n1 20.689
R11715 WE.n0 WE.t7 240.77
R11716 WE.n30 WE.t8 239.222
R11717 WE.n29 WE.t2 239.222
R11718 WE.n28 WE.t14 239.222
R11719 WE.n27 WE.t9 239.222
R11720 WE.n26 WE.t24 239.222
R11721 WE.n25 WE.t21 239.222
R11722 WE.n24 WE.t4 239.222
R11723 WE.n23 WE.t11 239.222
R11724 WE.n22 WE.t26 239.222
R11725 WE.n21 WE.t22 239.222
R11726 WE.n20 WE.t5 239.222
R11727 WE.n19 WE.t28 239.222
R11728 WE.n18 WE.t15 239.222
R11729 WE.n17 WE.t10 239.222
R11730 WE.n16 WE.t25 239.222
R11731 WE.n15 WE.t30 239.222
R11732 WE.n14 WE.t13 239.222
R11733 WE.n13 WE.t12 239.222
R11734 WE.n12 WE.t27 239.222
R11735 WE.n11 WE.t18 239.222
R11736 WE.n10 WE.t0 239.222
R11737 WE.n9 WE.t29 239.222
R11738 WE.n8 WE.t16 239.222
R11739 WE.n7 WE.t20 239.222
R11740 WE.n6 WE.t3 239.222
R11741 WE.n5 WE.t31 239.222
R11742 WE.n4 WE.t17 239.222
R11743 WE.n3 WE.t6 239.222
R11744 WE.n2 WE.t23 239.222
R11745 WE.n1 WE.t19 239.222
R11746 WE.n0 WE.t1 239.222
R11747 WE WE.n30 44.463
R11748 WE.n1 WE.n0 3.325
R11749 WE.n3 WE.n2 3.325
R11750 WE.n5 WE.n4 3.325
R11751 WE.n7 WE.n6 3.325
R11752 WE.n9 WE.n8 3.325
R11753 WE.n11 WE.n10 3.325
R11754 WE.n13 WE.n12 3.325
R11755 WE.n15 WE.n14 3.325
R11756 WE.n17 WE.n16 3.325
R11757 WE.n19 WE.n18 3.325
R11758 WE.n21 WE.n20 3.325
R11759 WE.n23 WE.n22 3.325
R11760 WE.n25 WE.n24 3.325
R11761 WE.n27 WE.n26 3.325
R11762 WE.n29 WE.n28 3.325
R11763 WE.n2 WE.n1 1.548
R11764 WE.n4 WE.n3 1.548
R11765 WE.n6 WE.n5 1.548
R11766 WE.n8 WE.n7 1.548
R11767 WE.n10 WE.n9 1.548
R11768 WE.n12 WE.n11 1.548
R11769 WE.n14 WE.n13 1.548
R11770 WE.n16 WE.n15 1.548
R11771 WE.n18 WE.n17 1.548
R11772 WE.n20 WE.n19 1.548
R11773 WE.n22 WE.n21 1.548
R11774 WE.n24 WE.n23 1.548
R11775 WE.n26 WE.n25 1.548
R11776 WE.n28 WE.n27 1.548
R11777 WE.n30 WE.n29 1.548
R11778 a_6133_n953.n25 a_6133_n953.t27 561.971
R11779 a_6133_n953.n0 a_6133_n953.t22 461.908
R11780 a_6133_n953.t7 a_6133_n953.n25 108.635
R11781 a_6133_n953.n0 a_6133_n953.t21 79.512
R11782 a_6133_n953.n24 a_6133_n953.t26 65.401
R11783 a_6133_n953.n23 a_6133_n953.t9 65.401
R11784 a_6133_n953.n22 a_6133_n953.t4 65.401
R11785 a_6133_n953.n21 a_6133_n953.t17 65.401
R11786 a_6133_n953.n20 a_6133_n953.t12 65.401
R11787 a_6133_n953.n19 a_6133_n953.t18 65.401
R11788 a_6133_n953.n18 a_6133_n953.t20 65.401
R11789 a_6133_n953.n17 a_6133_n953.t15 65.401
R11790 a_6133_n953.n16 a_6133_n953.t23 65.401
R11791 a_6133_n953.n15 a_6133_n953.t5 65.401
R11792 a_6133_n953.n14 a_6133_n953.t14 65.401
R11793 a_6133_n953.n13 a_6133_n953.t1 65.401
R11794 a_6133_n953.n12 a_6133_n953.t8 65.401
R11795 a_6133_n953.n11 a_6133_n953.t2 65.401
R11796 a_6133_n953.n10 a_6133_n953.t3 65.401
R11797 a_6133_n953.n9 a_6133_n953.t11 65.401
R11798 a_6133_n953.n8 a_6133_n953.t10 65.401
R11799 a_6133_n953.n7 a_6133_n953.t24 65.401
R11800 a_6133_n953.n6 a_6133_n953.t0 65.401
R11801 a_6133_n953.n5 a_6133_n953.t25 65.401
R11802 a_6133_n953.n4 a_6133_n953.t6 65.401
R11803 a_6133_n953.n3 a_6133_n953.t13 65.401
R11804 a_6133_n953.n2 a_6133_n953.t16 65.401
R11805 a_6133_n953.n1 a_6133_n953.t19 65.401
R11806 a_6133_n953.n1 a_6133_n953.n0 5.64
R11807 a_6133_n953.n25 a_6133_n953.n24 4.438
R11808 a_6133_n953.n23 a_6133_n953.n22 2.524
R11809 a_6133_n953.n3 a_6133_n953.n2 2.498
R11810 a_6133_n953.n17 a_6133_n953.n16 2.364
R11811 a_6133_n953.n9 a_6133_n953.n8 2.355
R11812 a_6133_n953.n2 a_6133_n953.n1 1.998
R11813 a_6133_n953.n4 a_6133_n953.n3 1.998
R11814 a_6133_n953.n5 a_6133_n953.n4 1.998
R11815 a_6133_n953.n6 a_6133_n953.n5 1.998
R11816 a_6133_n953.n7 a_6133_n953.n6 1.998
R11817 a_6133_n953.n8 a_6133_n953.n7 1.998
R11818 a_6133_n953.n10 a_6133_n953.n9 1.998
R11819 a_6133_n953.n11 a_6133_n953.n10 1.998
R11820 a_6133_n953.n12 a_6133_n953.n11 1.998
R11821 a_6133_n953.n13 a_6133_n953.n12 1.998
R11822 a_6133_n953.n14 a_6133_n953.n13 1.998
R11823 a_6133_n953.n15 a_6133_n953.n14 1.998
R11824 a_6133_n953.n16 a_6133_n953.n15 1.998
R11825 a_6133_n953.n18 a_6133_n953.n17 1.998
R11826 a_6133_n953.n19 a_6133_n953.n18 1.998
R11827 a_6133_n953.n20 a_6133_n953.n19 1.998
R11828 a_6133_n953.n21 a_6133_n953.n20 1.998
R11829 a_6133_n953.n22 a_6133_n953.n21 1.998
R11830 a_6133_n953.n24 a_6133_n953.n23 1.998
R11831 a_6203_n2086.t0 a_6203_n2086.t1 34.8
R11832 a_8997_n1053.n0 a_8997_n1053.t2 358.166
R11833 a_8997_n1053.t4 a_8997_n1053.t5 337.399
R11834 a_8997_n1053.t5 a_8997_n1053.t3 285.986
R11835 a_8997_n1053.n0 a_8997_n1053.t4 282.573
R11836 a_8997_n1053.n1 a_8997_n1053.t1 202.857
R11837 a_8997_n1053.n1 a_8997_n1053.n0 173.817
R11838 a_8997_n1053.n1 a_8997_n1053.t0 20.826
R11839 a_8997_n1053.n2 a_8997_n1053.n1 20.689
R11840 a_9367_n1053.t0 a_9367_n1053.t1 242.857
R11841 a_3247_3907.n0 a_3247_3907.t2 358.166
R11842 a_3247_3907.t4 a_3247_3907.t5 337.399
R11843 a_3247_3907.t5 a_3247_3907.t3 285.986
R11844 a_3247_3907.n0 a_3247_3907.t4 282.573
R11845 a_3247_3907.n1 a_3247_3907.t0 202.857
R11846 a_3247_3907.n1 a_3247_3907.n0 173.817
R11847 a_3247_3907.n1 a_3247_3907.t1 20.826
R11848 a_3247_3907.n2 a_3247_3907.n1 20.689
R11849 a_3258_n953.n25 a_3258_n953.t27 561.971
R11850 a_3258_n953.n0 a_3258_n953.t20 461.908
R11851 a_3258_n953.t5 a_3258_n953.n25 108.635
R11852 a_3258_n953.n0 a_3258_n953.t21 79.512
R11853 a_3258_n953.n24 a_3258_n953.t23 65.401
R11854 a_3258_n953.n23 a_3258_n953.t7 65.401
R11855 a_3258_n953.n22 a_3258_n953.t2 65.401
R11856 a_3258_n953.n21 a_3258_n953.t17 65.401
R11857 a_3258_n953.n20 a_3258_n953.t10 65.401
R11858 a_3258_n953.n19 a_3258_n953.t18 65.401
R11859 a_3258_n953.n18 a_3258_n953.t22 65.401
R11860 a_3258_n953.n17 a_3258_n953.t15 65.401
R11861 a_3258_n953.n16 a_3258_n953.t26 65.401
R11862 a_3258_n953.n15 a_3258_n953.t3 65.401
R11863 a_3258_n953.n14 a_3258_n953.t14 65.401
R11864 a_3258_n953.n13 a_3258_n953.t12 65.401
R11865 a_3258_n953.n12 a_3258_n953.t6 65.401
R11866 a_3258_n953.n11 a_3258_n953.t13 65.401
R11867 a_3258_n953.n10 a_3258_n953.t1 65.401
R11868 a_3258_n953.n9 a_3258_n953.t9 65.401
R11869 a_3258_n953.n8 a_3258_n953.t8 65.401
R11870 a_3258_n953.n7 a_3258_n953.t24 65.401
R11871 a_3258_n953.n6 a_3258_n953.t0 65.401
R11872 a_3258_n953.n5 a_3258_n953.t25 65.401
R11873 a_3258_n953.n4 a_3258_n953.t4 65.401
R11874 a_3258_n953.n3 a_3258_n953.t11 65.401
R11875 a_3258_n953.n2 a_3258_n953.t16 65.401
R11876 a_3258_n953.n1 a_3258_n953.t19 65.401
R11877 a_3258_n953.n1 a_3258_n953.n0 5.64
R11878 a_3258_n953.n25 a_3258_n953.n24 4.438
R11879 a_3258_n953.n23 a_3258_n953.n22 2.524
R11880 a_3258_n953.n3 a_3258_n953.n2 2.498
R11881 a_3258_n953.n17 a_3258_n953.n16 2.364
R11882 a_3258_n953.n9 a_3258_n953.n8 2.355
R11883 a_3258_n953.n2 a_3258_n953.n1 1.998
R11884 a_3258_n953.n4 a_3258_n953.n3 1.998
R11885 a_3258_n953.n5 a_3258_n953.n4 1.998
R11886 a_3258_n953.n6 a_3258_n953.n5 1.998
R11887 a_3258_n953.n7 a_3258_n953.n6 1.998
R11888 a_3258_n953.n8 a_3258_n953.n7 1.998
R11889 a_3258_n953.n10 a_3258_n953.n9 1.998
R11890 a_3258_n953.n11 a_3258_n953.n10 1.998
R11891 a_3258_n953.n12 a_3258_n953.n11 1.998
R11892 a_3258_n953.n13 a_3258_n953.n12 1.998
R11893 a_3258_n953.n14 a_3258_n953.n13 1.998
R11894 a_3258_n953.n15 a_3258_n953.n14 1.998
R11895 a_3258_n953.n16 a_3258_n953.n15 1.998
R11896 a_3258_n953.n18 a_3258_n953.n17 1.998
R11897 a_3258_n953.n19 a_3258_n953.n18 1.998
R11898 a_3258_n953.n20 a_3258_n953.n19 1.998
R11899 a_3258_n953.n21 a_3258_n953.n20 1.998
R11900 a_3258_n953.n22 a_3258_n953.n21 1.998
R11901 a_3258_n953.n24 a_3258_n953.n23 1.998
R11902 WWL[0].n0 WWL[0].t20 262.032
R11903 WWL[0].n29 WWL[0].t23 260.715
R11904 WWL[0].n27 WWL[0].t26 260.715
R11905 WWL[0].n25 WWL[0].t8 260.715
R11906 WWL[0].n23 WWL[0].t2 260.715
R11907 WWL[0].n21 WWL[0].t14 260.715
R11908 WWL[0].n19 WWL[0].t31 260.715
R11909 WWL[0].n17 WWL[0].t22 260.715
R11910 WWL[0].n15 WWL[0].t5 260.715
R11911 WWL[0].n13 WWL[0].t27 260.715
R11912 WWL[0].n11 WWL[0].t3 260.715
R11913 WWL[0].n9 WWL[0].t24 260.715
R11914 WWL[0].n7 WWL[0].t6 260.715
R11915 WWL[0].n5 WWL[0].t0 260.715
R11916 WWL[0].n3 WWL[0].t15 260.715
R11917 WWL[0].n1 WWL[0].t28 260.715
R11918 WWL[0].n30 WWL[0].t7 259.254
R11919 WWL[0].n28 WWL[0].t13 259.254
R11920 WWL[0].n26 WWL[0].t25 259.254
R11921 WWL[0].n24 WWL[0].t9 259.254
R11922 WWL[0].n22 WWL[0].t1 259.254
R11923 WWL[0].n20 WWL[0].t16 259.254
R11924 WWL[0].n18 WWL[0].t29 259.254
R11925 WWL[0].n16 WWL[0].t11 259.254
R11926 WWL[0].n14 WWL[0].t4 259.254
R11927 WWL[0].n12 WWL[0].t19 259.254
R11928 WWL[0].n10 WWL[0].t10 259.254
R11929 WWL[0].n8 WWL[0].t17 259.254
R11930 WWL[0].n6 WWL[0].t18 259.254
R11931 WWL[0].n4 WWL[0].t21 259.254
R11932 WWL[0].n2 WWL[0].t12 259.254
R11933 WWL[0].n0 WWL[0].t30 259.254
R11934 WWL[0] WWL[0].n30 44.647
R11935 WWL[0].n1 WWL[0].n0 3.576
R11936 WWL[0].n3 WWL[0].n2 3.576
R11937 WWL[0].n5 WWL[0].n4 3.576
R11938 WWL[0].n7 WWL[0].n6 3.576
R11939 WWL[0].n9 WWL[0].n8 3.576
R11940 WWL[0].n11 WWL[0].n10 3.576
R11941 WWL[0].n13 WWL[0].n12 3.576
R11942 WWL[0].n15 WWL[0].n14 3.576
R11943 WWL[0].n17 WWL[0].n16 3.576
R11944 WWL[0].n19 WWL[0].n18 3.576
R11945 WWL[0].n21 WWL[0].n20 3.576
R11946 WWL[0].n23 WWL[0].n22 3.576
R11947 WWL[0].n25 WWL[0].n24 3.576
R11948 WWL[0].n27 WWL[0].n26 3.576
R11949 WWL[0].n29 WWL[0].n28 3.576
R11950 WWL[0].n2 WWL[0].n1 1.317
R11951 WWL[0].n4 WWL[0].n3 1.317
R11952 WWL[0].n6 WWL[0].n5 1.317
R11953 WWL[0].n8 WWL[0].n7 1.317
R11954 WWL[0].n10 WWL[0].n9 1.317
R11955 WWL[0].n12 WWL[0].n11 1.317
R11956 WWL[0].n14 WWL[0].n13 1.317
R11957 WWL[0].n16 WWL[0].n15 1.317
R11958 WWL[0].n18 WWL[0].n17 1.317
R11959 WWL[0].n20 WWL[0].n19 1.317
R11960 WWL[0].n22 WWL[0].n21 1.317
R11961 WWL[0].n24 WWL[0].n23 1.317
R11962 WWL[0].n26 WWL[0].n25 1.317
R11963 WWL[0].n28 WWL[0].n27 1.317
R11964 WWL[0].n30 WWL[0].n29 1.317
R11965 a_7445_4887.n25 a_7445_4887.t27 561.971
R11966 a_7445_4887.n0 a_7445_4887.t22 449.944
R11967 a_7445_4887.t6 a_7445_4887.n25 108.636
R11968 a_7445_4887.n0 a_7445_4887.t21 74.821
R11969 a_7445_4887.n24 a_7445_4887.t26 63.519
R11970 a_7445_4887.n23 a_7445_4887.t8 63.519
R11971 a_7445_4887.n22 a_7445_4887.t2 63.519
R11972 a_7445_4887.n21 a_7445_4887.t18 63.519
R11973 a_7445_4887.n20 a_7445_4887.t11 63.519
R11974 a_7445_4887.n19 a_7445_4887.t19 63.519
R11975 a_7445_4887.n18 a_7445_4887.t24 63.519
R11976 a_7445_4887.n17 a_7445_4887.t16 63.519
R11977 a_7445_4887.n16 a_7445_4887.t23 63.519
R11978 a_7445_4887.n15 a_7445_4887.t3 63.519
R11979 a_7445_4887.n14 a_7445_4887.t15 63.519
R11980 a_7445_4887.n13 a_7445_4887.t0 63.519
R11981 a_7445_4887.n12 a_7445_4887.t7 63.519
R11982 a_7445_4887.n11 a_7445_4887.t13 63.519
R11983 a_7445_4887.n10 a_7445_4887.t5 63.519
R11984 a_7445_4887.n9 a_7445_4887.t10 63.519
R11985 a_7445_4887.n8 a_7445_4887.t9 63.519
R11986 a_7445_4887.n7 a_7445_4887.t25 63.519
R11987 a_7445_4887.n6 a_7445_4887.t1 63.519
R11988 a_7445_4887.n5 a_7445_4887.t14 63.519
R11989 a_7445_4887.n4 a_7445_4887.t4 63.519
R11990 a_7445_4887.n3 a_7445_4887.t12 63.519
R11991 a_7445_4887.n2 a_7445_4887.t17 63.519
R11992 a_7445_4887.n1 a_7445_4887.t20 63.519
R11993 a_7445_4887.n1 a_7445_4887.n0 8.619
R11994 a_7445_4887.n25 a_7445_4887.n24 2.946
R11995 a_7445_4887.n23 a_7445_4887.n22 2.524
R11996 a_7445_4887.n3 a_7445_4887.n2 2.498
R11997 a_7445_4887.n17 a_7445_4887.n16 2.364
R11998 a_7445_4887.n9 a_7445_4887.n8 2.355
R11999 a_7445_4887.n24 a_7445_4887.n23 1.998
R12000 a_7445_4887.n22 a_7445_4887.n21 1.998
R12001 a_7445_4887.n21 a_7445_4887.n20 1.998
R12002 a_7445_4887.n20 a_7445_4887.n19 1.998
R12003 a_7445_4887.n19 a_7445_4887.n18 1.998
R12004 a_7445_4887.n18 a_7445_4887.n17 1.998
R12005 a_7445_4887.n16 a_7445_4887.n15 1.998
R12006 a_7445_4887.n15 a_7445_4887.n14 1.998
R12007 a_7445_4887.n14 a_7445_4887.n13 1.998
R12008 a_7445_4887.n13 a_7445_4887.n12 1.998
R12009 a_7445_4887.n12 a_7445_4887.n11 1.998
R12010 a_7445_4887.n11 a_7445_4887.n10 1.998
R12011 a_7445_4887.n10 a_7445_4887.n9 1.998
R12012 a_7445_4887.n8 a_7445_4887.n7 1.998
R12013 a_7445_4887.n7 a_7445_4887.n6 1.998
R12014 a_7445_4887.n6 a_7445_4887.n5 1.998
R12015 a_7445_4887.n5 a_7445_4887.n4 1.998
R12016 a_7445_4887.n4 a_7445_4887.n3 1.998
R12017 a_7445_4887.n2 a_7445_4887.n1 1.998
R12018 a_7177_3651.n0 a_7177_3651.t2 362.857
R12019 a_7177_3651.t3 a_7177_3651.t4 337.399
R12020 a_7177_3651.t4 a_7177_3651.t5 298.839
R12021 a_7177_3651.n0 a_7177_3651.t3 280.405
R12022 a_7177_3651.n1 a_7177_3651.t0 200
R12023 a_7177_3651.n1 a_7177_3651.n0 172.311
R12024 a_7177_3651.n2 a_7177_3651.n1 24
R12025 a_7177_3651.n1 a_7177_3651.t1 21.212
R12026 a_4877_n286.n0 a_4877_n286.t0 362.857
R12027 a_4877_n286.t5 a_4877_n286.t4 337.399
R12028 a_4877_n286.t4 a_4877_n286.t3 298.839
R12029 a_4877_n286.n0 a_4877_n286.t5 280.405
R12030 a_4877_n286.n1 a_4877_n286.t2 200
R12031 a_4877_n286.n1 a_4877_n286.n0 172.311
R12032 a_4877_n286.n2 a_4877_n286.n1 24
R12033 a_4877_n286.n1 a_4877_n286.t1 21.212
R12034 a_4890_n271.t0 a_4890_n271.t1 242.857
R12035 a_7177_n286.n0 a_7177_n286.t1 362.857
R12036 a_7177_n286.t3 a_7177_n286.t4 337.399
R12037 a_7177_n286.t4 a_7177_n286.t5 298.839
R12038 a_7177_n286.n0 a_7177_n286.t3 280.405
R12039 a_7177_n286.n1 a_7177_n286.t0 200
R12040 a_7177_n286.n1 a_7177_n286.n0 172.311
R12041 a_7177_n286.n2 a_7177_n286.n1 24
R12042 a_7177_n286.n1 a_7177_n286.t2 21.212
R12043 a_7272_n271.n0 a_7272_n271.t1 358.166
R12044 a_7272_n271.t3 a_7272_n271.t5 337.399
R12045 a_7272_n271.t5 a_7272_n271.t4 285.986
R12046 a_7272_n271.n0 a_7272_n271.t3 282.573
R12047 a_7272_n271.n1 a_7272_n271.t2 202.857
R12048 a_7272_n271.n1 a_7272_n271.n0 173.817
R12049 a_7272_n271.n1 a_7272_n271.t0 20.826
R12050 a_7272_n271.n2 a_7272_n271.n1 20.689
R12051 a_2672_n512.n0 a_2672_n512.t2 358.166
R12052 a_2672_n512.t3 a_2672_n512.t4 337.399
R12053 a_2672_n512.t4 a_2672_n512.t5 285.986
R12054 a_2672_n512.n0 a_2672_n512.t3 282.573
R12055 a_2672_n512.n1 a_2672_n512.t0 202.857
R12056 a_2672_n512.n1 a_2672_n512.n0 173.817
R12057 a_2672_n512.n1 a_2672_n512.t1 20.826
R12058 a_2672_n512.n2 a_2672_n512.n1 20.689
R12059 a_2577_n527.n0 a_2577_n527.t2 362.857
R12060 a_2577_n527.t5 a_2577_n527.t3 337.399
R12061 a_2577_n527.t3 a_2577_n527.t4 298.839
R12062 a_2577_n527.n0 a_2577_n527.t5 280.405
R12063 a_2577_n527.n1 a_2577_n527.t0 200
R12064 a_2577_n527.n1 a_2577_n527.n0 172.311
R12065 a_2577_n527.n2 a_2577_n527.n1 24
R12066 a_2577_n527.n1 a_2577_n527.t1 21.212
R12067 a_8422_975.n0 a_8422_975.t1 358.166
R12068 a_8422_975.t4 a_8422_975.t3 337.399
R12069 a_8422_975.t3 a_8422_975.t5 285.986
R12070 a_8422_975.n0 a_8422_975.t4 282.573
R12071 a_8422_975.n1 a_8422_975.t2 202.857
R12072 a_8422_975.n1 a_8422_975.n0 173.817
R12073 a_8422_975.n1 a_8422_975.t0 20.826
R12074 a_8422_975.n2 a_8422_975.n1 20.689
R12075 a_8327_960.n0 a_8327_960.t1 362.857
R12076 a_8327_960.t4 a_8327_960.t3 337.399
R12077 a_8327_960.t3 a_8327_960.t5 298.839
R12078 a_8327_960.n0 a_8327_960.t4 280.405
R12079 a_8327_960.n1 a_8327_960.t2 200
R12080 a_8327_960.n1 a_8327_960.n0 172.311
R12081 a_8327_960.n2 a_8327_960.n1 24
R12082 a_8327_960.n1 a_8327_960.t0 21.212
R12083 a_3152_n1068.n0 a_3152_n1068.t0 362.857
R12084 a_3152_n1068.t3 a_3152_n1068.t4 337.399
R12085 a_3152_n1068.t4 a_3152_n1068.t5 298.839
R12086 a_3152_n1068.n0 a_3152_n1068.t3 280.405
R12087 a_3152_n1068.n1 a_3152_n1068.t2 200
R12088 a_3152_n1068.n1 a_3152_n1068.n0 172.311
R12089 a_3152_n1068.n2 a_3152_n1068.n1 24
R12090 a_3152_n1068.n1 a_3152_n1068.t1 21.212
R12091 a_3247_n1053.n0 a_3247_n1053.t1 358.166
R12092 a_3247_n1053.t4 a_3247_n1053.t5 337.399
R12093 a_3247_n1053.t5 a_3247_n1053.t3 285.986
R12094 a_3247_n1053.n0 a_3247_n1053.t4 282.573
R12095 a_3247_n1053.n1 a_3247_n1053.t2 202.857
R12096 a_3247_n1053.n1 a_3247_n1053.n0 173.817
R12097 a_3247_n1053.n1 a_3247_n1053.t0 20.826
R12098 a_3247_n1053.n2 a_3247_n1053.n1 20.689
R12099 a_2577_n1068.n0 a_2577_n1068.t0 362.857
R12100 a_2577_n1068.t5 a_2577_n1068.t3 337.399
R12101 a_2577_n1068.t3 a_2577_n1068.t4 298.839
R12102 a_2577_n1068.n0 a_2577_n1068.t5 280.405
R12103 a_2577_n1068.n1 a_2577_n1068.t2 200
R12104 a_2577_n1068.n1 a_2577_n1068.n0 172.311
R12105 a_2577_n1068.n2 a_2577_n1068.n1 24
R12106 a_2577_n1068.n1 a_2577_n1068.t1 21.212
R12107 a_2672_n1053.n0 a_2672_n1053.t1 358.166
R12108 a_2672_n1053.t5 a_2672_n1053.t3 337.399
R12109 a_2672_n1053.t3 a_2672_n1053.t4 285.986
R12110 a_2672_n1053.n0 a_2672_n1053.t5 282.573
R12111 a_2672_n1053.n1 a_2672_n1053.t2 202.857
R12112 a_2672_n1053.n1 a_2672_n1053.n0 173.817
R12113 a_2672_n1053.n1 a_2672_n1053.t0 20.826
R12114 a_2672_n1053.n2 a_2672_n1053.n1 20.689
R12115 a_3152_3651.n0 a_3152_3651.t2 362.857
R12116 a_3152_3651.t3 a_3152_3651.t4 337.399
R12117 a_3152_3651.t4 a_3152_3651.t5 298.839
R12118 a_3152_3651.n0 a_3152_3651.t3 280.405
R12119 a_3152_3651.n1 a_3152_3651.t0 200
R12120 a_3152_3651.n1 a_3152_3651.n0 172.311
R12121 a_3152_3651.n2 a_3152_3651.n1 24
R12122 a_3152_3651.n1 a_3152_3651.t1 21.212
R12123 a_8902_2647.n0 a_8902_2647.t1 362.857
R12124 a_8902_2647.t5 a_8902_2647.t4 337.399
R12125 a_8902_2647.t4 a_8902_2647.t3 298.839
R12126 a_8902_2647.n0 a_8902_2647.t5 280.405
R12127 a_8902_2647.n1 a_8902_2647.t0 200
R12128 a_8902_2647.n1 a_8902_2647.n0 172.311
R12129 a_8902_2647.n2 a_8902_2647.n1 24
R12130 a_8902_2647.n1 a_8902_2647.t2 21.212
R12131 a_8915_2662.t0 a_8915_2662.t1 242.857
R12132 a_4302_1683.n0 a_4302_1683.t2 362.857
R12133 a_4302_1683.t3 a_4302_1683.t5 337.399
R12134 a_4302_1683.t5 a_4302_1683.t4 298.839
R12135 a_4302_1683.n0 a_4302_1683.t3 280.405
R12136 a_4302_1683.n1 a_4302_1683.t0 200
R12137 a_4302_1683.n1 a_4302_1683.n0 172.311
R12138 a_4302_1683.n2 a_4302_1683.n1 24
R12139 a_4302_1683.n1 a_4302_1683.t1 21.212
R12140 SA_OUT[12].n1 SA_OUT[12].t3 661.027
R12141 SA_OUT[12].n1 SA_OUT[12].t4 392.255
R12142 SA_OUT[12].n2 SA_OUT[12].t2 223.716
R12143 SA_OUT[12].n0 SA_OUT[12].t0 153.977
R12144 SA_OUT[12].n2 SA_OUT[12].n1 143.764
R12145 SA_OUT[12].n0 SA_OUT[12].t1 59.86
R12146 SA_OUT[12] SA_OUT[12].n3 13.941
R12147 SA_OUT[12].n3 SA_OUT[12].n2 3.764
R12148 SA_OUT[12].n3 SA_OUT[12].n0 0.752
R12149 a_277_4430.n0 a_277_4430.t1 362.857
R12150 a_277_4430.t5 a_277_4430.t3 337.399
R12151 a_277_4430.t3 a_277_4430.t4 298.839
R12152 a_277_4430.n0 a_277_4430.t5 280.405
R12153 a_277_4430.n1 a_277_4430.t2 200
R12154 a_277_4430.n1 a_277_4430.n0 172.311
R12155 a_277_4430.n2 a_277_4430.n1 24
R12156 a_277_4430.n1 a_277_4430.t0 21.212
R12157 a_372_4445.n0 a_372_4445.t1 358.166
R12158 a_372_4445.t3 a_372_4445.t5 337.399
R12159 a_372_4445.t5 a_372_4445.t4 285.986
R12160 a_372_4445.n0 a_372_4445.t3 282.573
R12161 a_372_4445.n1 a_372_4445.t2 202.857
R12162 a_372_4445.n1 a_372_4445.n0 173.817
R12163 a_372_4445.n1 a_372_4445.t0 20.826
R12164 a_372_4445.n2 a_372_4445.n1 20.689
R12165 a_6027_2165.n0 a_6027_2165.t0 362.857
R12166 a_6027_2165.t4 a_6027_2165.t5 337.399
R12167 a_6027_2165.t5 a_6027_2165.t3 298.839
R12168 a_6027_2165.n0 a_6027_2165.t4 280.405
R12169 a_6027_2165.n1 a_6027_2165.t2 200
R12170 a_6027_2165.n1 a_6027_2165.n0 172.311
R12171 a_6027_2165.n2 a_6027_2165.n1 24
R12172 a_6027_2165.n1 a_6027_2165.t1 21.212
R12173 a_6040_2180.t0 a_6040_2180.t1 242.857
R12174 a_8422_1698.n0 a_8422_1698.t2 358.166
R12175 a_8422_1698.t5 a_8422_1698.t4 337.399
R12176 a_8422_1698.t4 a_8422_1698.t3 285.986
R12177 a_8422_1698.n0 a_8422_1698.t5 282.573
R12178 a_8422_1698.n1 a_8422_1698.t0 202.857
R12179 a_8422_1698.n1 a_8422_1698.n0 173.817
R12180 a_8422_1698.n1 a_8422_1698.t1 20.826
R12181 a_8422_1698.n2 a_8422_1698.n1 20.689
R12182 a_8792_1698.t0 a_8792_1698.t1 242.857
R12183 WWL[12].n0 WWL[12].t23 262.032
R12184 WWL[12].n29 WWL[12].t3 260.715
R12185 WWL[12].n27 WWL[12].t1 260.715
R12186 WWL[12].n25 WWL[12].t27 260.715
R12187 WWL[12].n23 WWL[12].t5 260.715
R12188 WWL[12].n21 WWL[12].t2 260.715
R12189 WWL[12].n19 WWL[12].t18 260.715
R12190 WWL[12].n17 WWL[12].t6 260.715
R12191 WWL[12].n15 WWL[12].t24 260.715
R12192 WWL[12].n13 WWL[12].t11 260.715
R12193 WWL[12].n11 WWL[12].t7 260.715
R12194 WWL[12].n9 WWL[12].t25 260.715
R12195 WWL[12].n7 WWL[12].t12 260.715
R12196 WWL[12].n5 WWL[12].t0 260.715
R12197 WWL[12].n3 WWL[12].t17 260.715
R12198 WWL[12].n1 WWL[12].t13 260.715
R12199 WWL[12].n30 WWL[12].t30 259.254
R12200 WWL[12].n28 WWL[12].t22 259.254
R12201 WWL[12].n26 WWL[12].t20 259.254
R12202 WWL[12].n24 WWL[12].t9 259.254
R12203 WWL[12].n22 WWL[12].t28 259.254
R12204 WWL[12].n20 WWL[12].t14 259.254
R12205 WWL[12].n18 WWL[12].t10 259.254
R12206 WWL[12].n16 WWL[12].t31 259.254
R12207 WWL[12].n14 WWL[12].t15 259.254
R12208 WWL[12].n12 WWL[12].t4 259.254
R12209 WWL[12].n10 WWL[12].t19 259.254
R12210 WWL[12].n8 WWL[12].t16 259.254
R12211 WWL[12].n6 WWL[12].t26 259.254
R12212 WWL[12].n4 WWL[12].t21 259.254
R12213 WWL[12].n2 WWL[12].t8 259.254
R12214 WWL[12].n0 WWL[12].t29 259.254
R12215 WWL[12] WWL[12].n30 44.647
R12216 WWL[12].n1 WWL[12].n0 3.576
R12217 WWL[12].n3 WWL[12].n2 3.576
R12218 WWL[12].n5 WWL[12].n4 3.576
R12219 WWL[12].n7 WWL[12].n6 3.576
R12220 WWL[12].n9 WWL[12].n8 3.576
R12221 WWL[12].n11 WWL[12].n10 3.576
R12222 WWL[12].n13 WWL[12].n12 3.576
R12223 WWL[12].n15 WWL[12].n14 3.576
R12224 WWL[12].n17 WWL[12].n16 3.576
R12225 WWL[12].n19 WWL[12].n18 3.576
R12226 WWL[12].n21 WWL[12].n20 3.576
R12227 WWL[12].n23 WWL[12].n22 3.576
R12228 WWL[12].n25 WWL[12].n24 3.576
R12229 WWL[12].n27 WWL[12].n26 3.576
R12230 WWL[12].n29 WWL[12].n28 3.576
R12231 WWL[12].n2 WWL[12].n1 1.317
R12232 WWL[12].n4 WWL[12].n3 1.317
R12233 WWL[12].n6 WWL[12].n5 1.317
R12234 WWL[12].n8 WWL[12].n7 1.317
R12235 WWL[12].n10 WWL[12].n9 1.317
R12236 WWL[12].n12 WWL[12].n11 1.317
R12237 WWL[12].n14 WWL[12].n13 1.317
R12238 WWL[12].n16 WWL[12].n15 1.317
R12239 WWL[12].n18 WWL[12].n17 1.317
R12240 WWL[12].n20 WWL[12].n19 1.317
R12241 WWL[12].n22 WWL[12].n21 1.317
R12242 WWL[12].n24 WWL[12].n23 1.317
R12243 WWL[12].n26 WWL[12].n25 1.317
R12244 WWL[12].n28 WWL[12].n27 1.317
R12245 WWL[12].n30 WWL[12].n29 1.317
R12246 a_7177_678.n0 a_7177_678.t1 362.857
R12247 a_7177_678.t4 a_7177_678.t3 337.399
R12248 a_7177_678.t3 a_7177_678.t5 298.839
R12249 a_7177_678.n0 a_7177_678.t4 280.405
R12250 a_7177_678.n1 a_7177_678.t0 200
R12251 a_7177_678.n1 a_7177_678.n0 172.311
R12252 a_7177_678.n2 a_7177_678.n1 24
R12253 a_7177_678.n1 a_7177_678.t2 21.212
R12254 a_3727_n827.n0 a_3727_n827.t1 362.857
R12255 a_3727_n827.t5 a_3727_n827.t3 337.399
R12256 a_3727_n827.t3 a_3727_n827.t4 298.839
R12257 a_3727_n827.n0 a_3727_n827.t5 280.405
R12258 a_3727_n827.n1 a_3727_n827.t0 200
R12259 a_3727_n827.n1 a_3727_n827.n0 172.311
R12260 a_3727_n827.n2 a_3727_n827.n1 24
R12261 a_3727_n827.n1 a_3727_n827.t2 21.212
R12262 a_3822_n812.n0 a_3822_n812.t1 358.166
R12263 a_3822_n812.t4 a_3822_n812.t3 337.399
R12264 a_3822_n812.t3 a_3822_n812.t5 285.986
R12265 a_3822_n812.n0 a_3822_n812.t4 282.573
R12266 a_3822_n812.n1 a_3822_n812.t2 202.857
R12267 a_3822_n812.n1 a_3822_n812.n0 173.817
R12268 a_3822_n812.n1 a_3822_n812.t0 20.826
R12269 a_3822_n812.n2 a_3822_n812.n1 20.689
R12270 a_7272_3666.n0 a_7272_3666.t1 358.166
R12271 a_7272_3666.t5 a_7272_3666.t4 337.399
R12272 a_7272_3666.t4 a_7272_3666.t3 285.986
R12273 a_7272_3666.n0 a_7272_3666.t5 282.573
R12274 a_7272_3666.n1 a_7272_3666.t2 202.857
R12275 a_7272_3666.n1 a_7272_3666.n0 173.817
R12276 a_7272_3666.n1 a_7272_3666.t0 20.826
R12277 a_7272_3666.n2 a_7272_3666.n1 20.689
R12278 a_7642_3666.t0 a_7642_3666.t1 242.857
R12279 a_8595_4887.n25 a_8595_4887.t27 561.971
R12280 a_8595_4887.n0 a_8595_4887.t21 449.944
R12281 a_8595_4887.t6 a_8595_4887.n25 108.636
R12282 a_8595_4887.n0 a_8595_4887.t22 74.821
R12283 a_8595_4887.n24 a_8595_4887.t25 63.519
R12284 a_8595_4887.n23 a_8595_4887.t8 63.519
R12285 a_8595_4887.n22 a_8595_4887.t2 63.519
R12286 a_8595_4887.n21 a_8595_4887.t18 63.519
R12287 a_8595_4887.n20 a_8595_4887.t11 63.519
R12288 a_8595_4887.n19 a_8595_4887.t19 63.519
R12289 a_8595_4887.n18 a_8595_4887.t23 63.519
R12290 a_8595_4887.n17 a_8595_4887.t5 63.519
R12291 a_8595_4887.n16 a_8595_4887.t26 63.519
R12292 a_8595_4887.n15 a_8595_4887.t3 63.519
R12293 a_8595_4887.n14 a_8595_4887.t16 63.519
R12294 a_8595_4887.n13 a_8595_4887.t12 63.519
R12295 a_8595_4887.n12 a_8595_4887.t7 63.519
R12296 a_8595_4887.n11 a_8595_4887.t14 63.519
R12297 a_8595_4887.n10 a_8595_4887.t1 63.519
R12298 a_8595_4887.n9 a_8595_4887.t10 63.519
R12299 a_8595_4887.n8 a_8595_4887.t9 63.519
R12300 a_8595_4887.n7 a_8595_4887.t24 63.519
R12301 a_8595_4887.n6 a_8595_4887.t0 63.519
R12302 a_8595_4887.n5 a_8595_4887.t15 63.519
R12303 a_8595_4887.n4 a_8595_4887.t4 63.519
R12304 a_8595_4887.n3 a_8595_4887.t13 63.519
R12305 a_8595_4887.n2 a_8595_4887.t17 63.519
R12306 a_8595_4887.n1 a_8595_4887.t20 63.519
R12307 a_8595_4887.n1 a_8595_4887.n0 8.619
R12308 a_8595_4887.n25 a_8595_4887.n24 2.946
R12309 a_8595_4887.n23 a_8595_4887.n22 2.524
R12310 a_8595_4887.n3 a_8595_4887.n2 2.498
R12311 a_8595_4887.n17 a_8595_4887.n16 2.364
R12312 a_8595_4887.n9 a_8595_4887.n8 2.355
R12313 a_8595_4887.n24 a_8595_4887.n23 1.998
R12314 a_8595_4887.n22 a_8595_4887.n21 1.998
R12315 a_8595_4887.n21 a_8595_4887.n20 1.998
R12316 a_8595_4887.n20 a_8595_4887.n19 1.998
R12317 a_8595_4887.n19 a_8595_4887.n18 1.998
R12318 a_8595_4887.n18 a_8595_4887.n17 1.998
R12319 a_8595_4887.n16 a_8595_4887.n15 1.998
R12320 a_8595_4887.n15 a_8595_4887.n14 1.998
R12321 a_8595_4887.n14 a_8595_4887.n13 1.998
R12322 a_8595_4887.n13 a_8595_4887.n12 1.998
R12323 a_8595_4887.n12 a_8595_4887.n11 1.998
R12324 a_8595_4887.n11 a_8595_4887.n10 1.998
R12325 a_8595_4887.n10 a_8595_4887.n9 1.998
R12326 a_8595_4887.n8 a_8595_4887.n7 1.998
R12327 a_8595_4887.n7 a_8595_4887.n6 1.998
R12328 a_8595_4887.n6 a_8595_4887.n5 1.998
R12329 a_8595_4887.n5 a_8595_4887.n4 1.998
R12330 a_8595_4887.n4 a_8595_4887.n3 1.998
R12331 a_8595_4887.n2 a_8595_4887.n1 1.998
R12332 a_8327_1924.n0 a_8327_1924.t2 362.857
R12333 a_8327_1924.t3 a_8327_1924.t4 337.399
R12334 a_8327_1924.t4 a_8327_1924.t5 298.839
R12335 a_8327_1924.n0 a_8327_1924.t3 280.405
R12336 a_8327_1924.n1 a_8327_1924.t0 200
R12337 a_8327_1924.n1 a_8327_1924.n0 172.311
R12338 a_8327_1924.n2 a_8327_1924.n1 24
R12339 a_8327_1924.n1 a_8327_1924.t1 21.212
R12340 a_4302_n827.n0 a_4302_n827.t1 362.857
R12341 a_4302_n827.t3 a_4302_n827.t5 337.399
R12342 a_4302_n827.t5 a_4302_n827.t4 298.839
R12343 a_4302_n827.n0 a_4302_n827.t3 280.405
R12344 a_4302_n827.n1 a_4302_n827.t2 200
R12345 a_4302_n827.n1 a_4302_n827.n0 172.311
R12346 a_4302_n827.n2 a_4302_n827.n1 24
R12347 a_4302_n827.n1 a_4302_n827.t0 21.212
R12348 a_7752_3410.n0 a_7752_3410.t1 362.857
R12349 a_7752_3410.t3 a_7752_3410.t4 337.399
R12350 a_7752_3410.t4 a_7752_3410.t5 298.839
R12351 a_7752_3410.n0 a_7752_3410.t3 280.405
R12352 a_7752_3410.n1 a_7752_3410.t0 200
R12353 a_7752_3410.n1 a_7752_3410.n0 172.311
R12354 a_7752_3410.n2 a_7752_3410.n1 24
R12355 a_7752_3410.n1 a_7752_3410.t2 21.212
R12356 RWL[3].n0 RWL[3].t14 154.243
R12357 RWL[3].n14 RWL[3].t4 149.249
R12358 RWL[3].n13 RWL[3].t9 149.249
R12359 RWL[3].n12 RWL[3].t0 149.249
R12360 RWL[3].n11 RWL[3].t5 149.249
R12361 RWL[3].n10 RWL[3].t2 149.249
R12362 RWL[3].n9 RWL[3].t10 149.249
R12363 RWL[3].n8 RWL[3].t1 149.249
R12364 RWL[3].n7 RWL[3].t7 149.249
R12365 RWL[3].n6 RWL[3].t3 149.249
R12366 RWL[3].n5 RWL[3].t13 149.249
R12367 RWL[3].n4 RWL[3].t6 149.249
R12368 RWL[3].n3 RWL[3].t11 149.249
R12369 RWL[3].n2 RWL[3].t12 149.249
R12370 RWL[3].n1 RWL[3].t15 149.249
R12371 RWL[3].n0 RWL[3].t8 149.249
R12372 RWL[3] RWL[3].n14 42.872
R12373 RWL[3].n1 RWL[3].n0 4.994
R12374 RWL[3].n2 RWL[3].n1 4.994
R12375 RWL[3].n3 RWL[3].n2 4.994
R12376 RWL[3].n4 RWL[3].n3 4.994
R12377 RWL[3].n5 RWL[3].n4 4.994
R12378 RWL[3].n6 RWL[3].n5 4.994
R12379 RWL[3].n7 RWL[3].n6 4.994
R12380 RWL[3].n8 RWL[3].n7 4.994
R12381 RWL[3].n9 RWL[3].n8 4.994
R12382 RWL[3].n10 RWL[3].n9 4.994
R12383 RWL[3].n11 RWL[3].n10 4.994
R12384 RWL[3].n12 RWL[3].n11 4.994
R12385 RWL[3].n13 RWL[3].n12 4.994
R12386 RWL[3].n14 RWL[3].n13 4.994
R12387 a_1440_2943.t0 a_1440_2943.t1 242.857
R12388 a_1440_n953.t37 a_1440_n953.n46 176.385
R12389 a_1440_n953.n22 a_1440_n953.t9 67.378
R12390 a_1440_n953.n0 a_1440_n953.t15 66.92
R12391 a_1440_n953.n1 a_1440_n953.t5 66.92
R12392 a_1440_n953.n2 a_1440_n953.t8 66.92
R12393 a_1440_n953.n3 a_1440_n953.t11 66.92
R12394 a_1440_n953.n4 a_1440_n953.t1 66.92
R12395 a_1440_n953.n5 a_1440_n953.t48 66.92
R12396 a_1440_n953.n6 a_1440_n953.t39 66.92
R12397 a_1440_n953.n7 a_1440_n953.t46 66.92
R12398 a_1440_n953.n8 a_1440_n953.t23 66.92
R12399 a_1440_n953.n9 a_1440_n953.t30 66.92
R12400 a_1440_n953.n10 a_1440_n953.t19 66.92
R12401 a_1440_n953.n11 a_1440_n953.t33 66.92
R12402 a_1440_n953.n12 a_1440_n953.t27 66.92
R12403 a_1440_n953.n13 a_1440_n953.t42 66.92
R12404 a_1440_n953.n14 a_1440_n953.t47 66.92
R12405 a_1440_n953.n15 a_1440_n953.t45 66.92
R12406 a_1440_n953.n16 a_1440_n953.t18 66.92
R12407 a_1440_n953.n17 a_1440_n953.t24 66.92
R12408 a_1440_n953.n18 a_1440_n953.t22 66.92
R12409 a_1440_n953.n19 a_1440_n953.t25 66.92
R12410 a_1440_n953.n20 a_1440_n953.t7 66.92
R12411 a_1440_n953.n21 a_1440_n953.t6 66.92
R12412 a_1440_n953.n22 a_1440_n953.t14 66.92
R12413 a_1440_n953.n23 a_1440_n953.t16 65.518
R12414 a_1440_n953.n45 a_1440_n953.t3 63.519
R12415 a_1440_n953.n44 a_1440_n953.t12 63.519
R12416 a_1440_n953.n43 a_1440_n953.t17 63.519
R12417 a_1440_n953.n42 a_1440_n953.t4 63.519
R12418 a_1440_n953.n41 a_1440_n953.t32 63.519
R12419 a_1440_n953.n40 a_1440_n953.t38 63.519
R12420 a_1440_n953.n39 a_1440_n953.t21 63.519
R12421 a_1440_n953.n38 a_1440_n953.t20 63.519
R12422 a_1440_n953.n37 a_1440_n953.t44 63.519
R12423 a_1440_n953.n36 a_1440_n953.t36 63.519
R12424 a_1440_n953.n35 a_1440_n953.t31 63.519
R12425 a_1440_n953.n34 a_1440_n953.t29 63.519
R12426 a_1440_n953.n33 a_1440_n953.t0 63.519
R12427 a_1440_n953.n32 a_1440_n953.t40 63.519
R12428 a_1440_n953.n31 a_1440_n953.t41 63.519
R12429 a_1440_n953.n30 a_1440_n953.t35 63.519
R12430 a_1440_n953.n29 a_1440_n953.t34 63.519
R12431 a_1440_n953.n28 a_1440_n953.t43 63.519
R12432 a_1440_n953.n27 a_1440_n953.t28 63.519
R12433 a_1440_n953.n26 a_1440_n953.t26 63.519
R12434 a_1440_n953.n25 a_1440_n953.t13 63.519
R12435 a_1440_n953.n24 a_1440_n953.t10 63.519
R12436 a_1440_n953.n23 a_1440_n953.t2 63.519
R12437 a_1440_n953.n46 a_1440_n953.n0 19.599
R12438 a_1440_n953.n46 a_1440_n953.n45 15.67
R12439 a_1440_n953.n44 a_1440_n953.n43 2.524
R12440 a_1440_n953.n24 a_1440_n953.n23 2.498
R12441 a_1440_n953.n21 a_1440_n953.n22 2.495
R12442 a_1440_n953.n1 a_1440_n953.n2 2.459
R12443 a_1440_n953.n38 a_1440_n953.n37 2.364
R12444 a_1440_n953.n30 a_1440_n953.n29 2.355
R12445 a_1440_n953.n7 a_1440_n953.n8 2.299
R12446 a_1440_n953.n15 a_1440_n953.n16 2.29
R12447 a_1440_n953.n16 a_1440_n953.n17 2.057
R12448 a_1440_n953.n8 a_1440_n953.n9 2.057
R12449 a_1440_n953.n2 a_1440_n953.n3 2.057
R12450 a_1440_n953.n0 a_1440_n953.n1 2.057
R12451 a_1440_n953.n45 a_1440_n953.n44 1.998
R12452 a_1440_n953.n43 a_1440_n953.n42 1.998
R12453 a_1440_n953.n42 a_1440_n953.n41 1.998
R12454 a_1440_n953.n41 a_1440_n953.n40 1.998
R12455 a_1440_n953.n40 a_1440_n953.n39 1.998
R12456 a_1440_n953.n39 a_1440_n953.n38 1.998
R12457 a_1440_n953.n37 a_1440_n953.n36 1.998
R12458 a_1440_n953.n36 a_1440_n953.n35 1.998
R12459 a_1440_n953.n35 a_1440_n953.n34 1.998
R12460 a_1440_n953.n34 a_1440_n953.n33 1.998
R12461 a_1440_n953.n33 a_1440_n953.n32 1.998
R12462 a_1440_n953.n32 a_1440_n953.n31 1.998
R12463 a_1440_n953.n31 a_1440_n953.n30 1.998
R12464 a_1440_n953.n29 a_1440_n953.n28 1.998
R12465 a_1440_n953.n28 a_1440_n953.n27 1.998
R12466 a_1440_n953.n27 a_1440_n953.n26 1.998
R12467 a_1440_n953.n26 a_1440_n953.n25 1.998
R12468 a_1440_n953.n25 a_1440_n953.n24 1.998
R12469 a_1440_n953.n20 a_1440_n953.n21 1.995
R12470 a_1440_n953.n19 a_1440_n953.n20 1.995
R12471 a_1440_n953.n18 a_1440_n953.n19 1.995
R12472 a_1440_n953.n17 a_1440_n953.n18 1.995
R12473 a_1440_n953.n14 a_1440_n953.n15 1.995
R12474 a_1440_n953.n13 a_1440_n953.n14 1.995
R12475 a_1440_n953.n12 a_1440_n953.n13 1.995
R12476 a_1440_n953.n11 a_1440_n953.n12 1.995
R12477 a_1440_n953.n10 a_1440_n953.n11 1.995
R12478 a_1440_n953.n9 a_1440_n953.n10 1.995
R12479 a_1440_n953.n6 a_1440_n953.n7 1.995
R12480 a_1440_n953.n5 a_1440_n953.n6 1.995
R12481 a_1440_n953.n4 a_1440_n953.n5 1.995
R12482 a_1440_n953.n3 a_1440_n953.n4 1.995
R12483 WWL[9].n0 WWL[9].t0 262.032
R12484 WWL[9].n29 WWL[9].t3 260.715
R12485 WWL[9].n27 WWL[9].t6 260.715
R12486 WWL[9].n25 WWL[9].t20 260.715
R12487 WWL[9].n23 WWL[9].t14 260.715
R12488 WWL[9].n21 WWL[9].t26 260.715
R12489 WWL[9].n19 WWL[9].t11 260.715
R12490 WWL[9].n17 WWL[9].t2 260.715
R12491 WWL[9].n15 WWL[9].t17 260.715
R12492 WWL[9].n13 WWL[9].t7 260.715
R12493 WWL[9].n11 WWL[9].t15 260.715
R12494 WWL[9].n9 WWL[9].t4 260.715
R12495 WWL[9].n7 WWL[9].t18 260.715
R12496 WWL[9].n5 WWL[9].t12 260.715
R12497 WWL[9].n3 WWL[9].t27 260.715
R12498 WWL[9].n1 WWL[9].t8 260.715
R12499 WWL[9].n30 WWL[9].t19 259.254
R12500 WWL[9].n28 WWL[9].t25 259.254
R12501 WWL[9].n26 WWL[9].t5 259.254
R12502 WWL[9].n24 WWL[9].t21 259.254
R12503 WWL[9].n22 WWL[9].t13 259.254
R12504 WWL[9].n20 WWL[9].t28 259.254
R12505 WWL[9].n18 WWL[9].t9 259.254
R12506 WWL[9].n16 WWL[9].t23 259.254
R12507 WWL[9].n14 WWL[9].t16 259.254
R12508 WWL[9].n12 WWL[9].t31 259.254
R12509 WWL[9].n10 WWL[9].t22 259.254
R12510 WWL[9].n8 WWL[9].t29 259.254
R12511 WWL[9].n6 WWL[9].t30 259.254
R12512 WWL[9].n4 WWL[9].t1 259.254
R12513 WWL[9].n2 WWL[9].t24 259.254
R12514 WWL[9].n0 WWL[9].t10 259.254
R12515 WWL[9] WWL[9].n30 44.647
R12516 WWL[9].n1 WWL[9].n0 3.576
R12517 WWL[9].n3 WWL[9].n2 3.576
R12518 WWL[9].n5 WWL[9].n4 3.576
R12519 WWL[9].n7 WWL[9].n6 3.576
R12520 WWL[9].n9 WWL[9].n8 3.576
R12521 WWL[9].n11 WWL[9].n10 3.576
R12522 WWL[9].n13 WWL[9].n12 3.576
R12523 WWL[9].n15 WWL[9].n14 3.576
R12524 WWL[9].n17 WWL[9].n16 3.576
R12525 WWL[9].n19 WWL[9].n18 3.576
R12526 WWL[9].n21 WWL[9].n20 3.576
R12527 WWL[9].n23 WWL[9].n22 3.576
R12528 WWL[9].n25 WWL[9].n24 3.576
R12529 WWL[9].n27 WWL[9].n26 3.576
R12530 WWL[9].n29 WWL[9].n28 3.576
R12531 WWL[9].n2 WWL[9].n1 1.317
R12532 WWL[9].n4 WWL[9].n3 1.317
R12533 WWL[9].n6 WWL[9].n5 1.317
R12534 WWL[9].n8 WWL[9].n7 1.317
R12535 WWL[9].n10 WWL[9].n9 1.317
R12536 WWL[9].n12 WWL[9].n11 1.317
R12537 WWL[9].n14 WWL[9].n13 1.317
R12538 WWL[9].n16 WWL[9].n15 1.317
R12539 WWL[9].n18 WWL[9].n17 1.317
R12540 WWL[9].n20 WWL[9].n19 1.317
R12541 WWL[9].n22 WWL[9].n21 1.317
R12542 WWL[9].n24 WWL[9].n23 1.317
R12543 WWL[9].n26 WWL[9].n25 1.317
R12544 WWL[9].n28 WWL[9].n27 1.317
R12545 WWL[9].n30 WWL[9].n29 1.317
R12546 a_9170_4887.n25 a_9170_4887.t27 561.971
R12547 a_9170_4887.n0 a_9170_4887.t23 449.944
R12548 a_9170_4887.t7 a_9170_4887.n25 108.636
R12549 a_9170_4887.n0 a_9170_4887.t22 74.821
R12550 a_9170_4887.n24 a_9170_4887.t25 63.519
R12551 a_9170_4887.n23 a_9170_4887.t9 63.519
R12552 a_9170_4887.n22 a_9170_4887.t3 63.519
R12553 a_9170_4887.n21 a_9170_4887.t18 63.519
R12554 a_9170_4887.n20 a_9170_4887.t14 63.519
R12555 a_9170_4887.n19 a_9170_4887.t19 63.519
R12556 a_9170_4887.n18 a_9170_4887.t21 63.519
R12557 a_9170_4887.n17 a_9170_4887.t6 63.519
R12558 a_9170_4887.n16 a_9170_4887.t26 63.519
R12559 a_9170_4887.n15 a_9170_4887.t4 63.519
R12560 a_9170_4887.n14 a_9170_4887.t11 63.519
R12561 a_9170_4887.n13 a_9170_4887.t1 63.519
R12562 a_9170_4887.n12 a_9170_4887.t8 63.519
R12563 a_9170_4887.n11 a_9170_4887.t15 63.519
R12564 a_9170_4887.n10 a_9170_4887.t2 63.519
R12565 a_9170_4887.n9 a_9170_4887.t12 63.519
R12566 a_9170_4887.n8 a_9170_4887.t10 63.519
R12567 a_9170_4887.n7 a_9170_4887.t24 63.519
R12568 a_9170_4887.n6 a_9170_4887.t0 63.519
R12569 a_9170_4887.n5 a_9170_4887.t16 63.519
R12570 a_9170_4887.n4 a_9170_4887.t5 63.519
R12571 a_9170_4887.n3 a_9170_4887.t13 63.519
R12572 a_9170_4887.n2 a_9170_4887.t17 63.519
R12573 a_9170_4887.n1 a_9170_4887.t20 63.519
R12574 a_9170_4887.n1 a_9170_4887.n0 8.619
R12575 a_9170_4887.n25 a_9170_4887.n24 2.946
R12576 a_9170_4887.n23 a_9170_4887.n22 2.524
R12577 a_9170_4887.n3 a_9170_4887.n2 2.498
R12578 a_9170_4887.n17 a_9170_4887.n16 2.364
R12579 a_9170_4887.n9 a_9170_4887.n8 2.355
R12580 a_9170_4887.n24 a_9170_4887.n23 1.998
R12581 a_9170_4887.n22 a_9170_4887.n21 1.998
R12582 a_9170_4887.n21 a_9170_4887.n20 1.998
R12583 a_9170_4887.n20 a_9170_4887.n19 1.998
R12584 a_9170_4887.n19 a_9170_4887.n18 1.998
R12585 a_9170_4887.n18 a_9170_4887.n17 1.998
R12586 a_9170_4887.n16 a_9170_4887.n15 1.998
R12587 a_9170_4887.n15 a_9170_4887.n14 1.998
R12588 a_9170_4887.n14 a_9170_4887.n13 1.998
R12589 a_9170_4887.n13 a_9170_4887.n12 1.998
R12590 a_9170_4887.n12 a_9170_4887.n11 1.998
R12591 a_9170_4887.n11 a_9170_4887.n10 1.998
R12592 a_9170_4887.n10 a_9170_4887.n9 1.998
R12593 a_9170_4887.n8 a_9170_4887.n7 1.998
R12594 a_9170_4887.n7 a_9170_4887.n6 1.998
R12595 a_9170_4887.n6 a_9170_4887.n5 1.998
R12596 a_9170_4887.n5 a_9170_4887.n4 1.998
R12597 a_9170_4887.n4 a_9170_4887.n3 1.998
R12598 a_9170_4887.n2 a_9170_4887.n1 1.998
R12599 a_8902_1442.n0 a_8902_1442.t1 362.857
R12600 a_8902_1442.t4 a_8902_1442.t3 337.399
R12601 a_8902_1442.t3 a_8902_1442.t5 298.839
R12602 a_8902_1442.n0 a_8902_1442.t4 280.405
R12603 a_8902_1442.n1 a_8902_1442.t0 200
R12604 a_8902_1442.n1 a_8902_1442.n0 172.311
R12605 a_8902_1442.n2 a_8902_1442.n1 24
R12606 a_8902_1442.n1 a_8902_1442.t2 21.212
R12607 WWL[14].n0 WWL[14].t1 262.032
R12608 WWL[14].n29 WWL[14].t13 260.715
R12609 WWL[14].n27 WWL[14].t11 260.715
R12610 WWL[14].n25 WWL[14].t5 260.715
R12611 WWL[14].n23 WWL[14].t15 260.715
R12612 WWL[14].n21 WWL[14].t12 260.715
R12613 WWL[14].n19 WWL[14].t28 260.715
R12614 WWL[14].n17 WWL[14].t16 260.715
R12615 WWL[14].n15 WWL[14].t2 260.715
R12616 WWL[14].n13 WWL[14].t21 260.715
R12617 WWL[14].n11 WWL[14].t17 260.715
R12618 WWL[14].n9 WWL[14].t3 260.715
R12619 WWL[14].n7 WWL[14].t22 260.715
R12620 WWL[14].n5 WWL[14].t10 260.715
R12621 WWL[14].n3 WWL[14].t27 260.715
R12622 WWL[14].n1 WWL[14].t23 260.715
R12623 WWL[14].n30 WWL[14].t8 259.254
R12624 WWL[14].n28 WWL[14].t0 259.254
R12625 WWL[14].n26 WWL[14].t30 259.254
R12626 WWL[14].n24 WWL[14].t19 259.254
R12627 WWL[14].n22 WWL[14].t6 259.254
R12628 WWL[14].n20 WWL[14].t24 259.254
R12629 WWL[14].n18 WWL[14].t20 259.254
R12630 WWL[14].n16 WWL[14].t9 259.254
R12631 WWL[14].n14 WWL[14].t25 259.254
R12632 WWL[14].n12 WWL[14].t14 259.254
R12633 WWL[14].n10 WWL[14].t29 259.254
R12634 WWL[14].n8 WWL[14].t26 259.254
R12635 WWL[14].n6 WWL[14].t4 259.254
R12636 WWL[14].n4 WWL[14].t31 259.254
R12637 WWL[14].n2 WWL[14].t18 259.254
R12638 WWL[14].n0 WWL[14].t7 259.254
R12639 WWL[14] WWL[14].n30 44.647
R12640 WWL[14].n1 WWL[14].n0 3.576
R12641 WWL[14].n3 WWL[14].n2 3.576
R12642 WWL[14].n5 WWL[14].n4 3.576
R12643 WWL[14].n7 WWL[14].n6 3.576
R12644 WWL[14].n9 WWL[14].n8 3.576
R12645 WWL[14].n11 WWL[14].n10 3.576
R12646 WWL[14].n13 WWL[14].n12 3.576
R12647 WWL[14].n15 WWL[14].n14 3.576
R12648 WWL[14].n17 WWL[14].n16 3.576
R12649 WWL[14].n19 WWL[14].n18 3.576
R12650 WWL[14].n21 WWL[14].n20 3.576
R12651 WWL[14].n23 WWL[14].n22 3.576
R12652 WWL[14].n25 WWL[14].n24 3.576
R12653 WWL[14].n27 WWL[14].n26 3.576
R12654 WWL[14].n29 WWL[14].n28 3.576
R12655 WWL[14].n2 WWL[14].n1 1.317
R12656 WWL[14].n4 WWL[14].n3 1.317
R12657 WWL[14].n6 WWL[14].n5 1.317
R12658 WWL[14].n8 WWL[14].n7 1.317
R12659 WWL[14].n10 WWL[14].n9 1.317
R12660 WWL[14].n12 WWL[14].n11 1.317
R12661 WWL[14].n14 WWL[14].n13 1.317
R12662 WWL[14].n16 WWL[14].n15 1.317
R12663 WWL[14].n18 WWL[14].n17 1.317
R12664 WWL[14].n20 WWL[14].n19 1.317
R12665 WWL[14].n22 WWL[14].n21 1.317
R12666 WWL[14].n24 WWL[14].n23 1.317
R12667 WWL[14].n26 WWL[14].n25 1.317
R12668 WWL[14].n28 WWL[14].n27 1.317
R12669 WWL[14].n30 WWL[14].n29 1.317
R12670 a_947_211.n0 a_947_211.t1 358.166
R12671 a_947_211.t4 a_947_211.t3 337.399
R12672 a_947_211.t3 a_947_211.t5 285.986
R12673 a_947_211.n0 a_947_211.t4 282.573
R12674 a_947_211.n1 a_947_211.t2 202.857
R12675 a_947_211.n1 a_947_211.n0 173.817
R12676 a_947_211.n1 a_947_211.t0 20.826
R12677 a_947_211.n2 a_947_211.n1 20.689
R12678 a_958_n953.n25 a_958_n953.t27 561.971
R12679 a_958_n953.n0 a_958_n953.t22 461.908
R12680 a_958_n953.t7 a_958_n953.n25 108.635
R12681 a_958_n953.n0 a_958_n953.t23 79.512
R12682 a_958_n953.n24 a_958_n953.t24 65.401
R12683 a_958_n953.n23 a_958_n953.t10 65.401
R12684 a_958_n953.n22 a_958_n953.t3 65.401
R12685 a_958_n953.n21 a_958_n953.t19 65.401
R12686 a_958_n953.n20 a_958_n953.t15 65.401
R12687 a_958_n953.n19 a_958_n953.t9 65.401
R12688 a_958_n953.n18 a_958_n953.t21 65.401
R12689 a_958_n953.n17 a_958_n953.t6 65.401
R12690 a_958_n953.n16 a_958_n953.t26 65.401
R12691 a_958_n953.n15 a_958_n953.t4 65.401
R12692 a_958_n953.n14 a_958_n953.t12 65.401
R12693 a_958_n953.n13 a_958_n953.t1 65.401
R12694 a_958_n953.n12 a_958_n953.t8 65.401
R12695 a_958_n953.n11 a_958_n953.t16 65.401
R12696 a_958_n953.n10 a_958_n953.t2 65.401
R12697 a_958_n953.n9 a_958_n953.t13 65.401
R12698 a_958_n953.n8 a_958_n953.t11 65.401
R12699 a_958_n953.n7 a_958_n953.t25 65.401
R12700 a_958_n953.n6 a_958_n953.t0 65.401
R12701 a_958_n953.n5 a_958_n953.t17 65.401
R12702 a_958_n953.n4 a_958_n953.t5 65.401
R12703 a_958_n953.n3 a_958_n953.t14 65.401
R12704 a_958_n953.n2 a_958_n953.t18 65.401
R12705 a_958_n953.n1 a_958_n953.t20 65.401
R12706 a_958_n953.n1 a_958_n953.n0 5.64
R12707 a_958_n953.n25 a_958_n953.n24 4.438
R12708 a_958_n953.n23 a_958_n953.n22 2.524
R12709 a_958_n953.n3 a_958_n953.n2 2.498
R12710 a_958_n953.n17 a_958_n953.n16 2.364
R12711 a_958_n953.n9 a_958_n953.n8 2.355
R12712 a_958_n953.n2 a_958_n953.n1 1.998
R12713 a_958_n953.n4 a_958_n953.n3 1.998
R12714 a_958_n953.n5 a_958_n953.n4 1.998
R12715 a_958_n953.n6 a_958_n953.n5 1.998
R12716 a_958_n953.n7 a_958_n953.n6 1.998
R12717 a_958_n953.n8 a_958_n953.n7 1.998
R12718 a_958_n953.n10 a_958_n953.n9 1.998
R12719 a_958_n953.n11 a_958_n953.n10 1.998
R12720 a_958_n953.n12 a_958_n953.n11 1.998
R12721 a_958_n953.n13 a_958_n953.n12 1.998
R12722 a_958_n953.n14 a_958_n953.n13 1.998
R12723 a_958_n953.n15 a_958_n953.n14 1.998
R12724 a_958_n953.n16 a_958_n953.n15 1.998
R12725 a_958_n953.n18 a_958_n953.n17 1.998
R12726 a_958_n953.n19 a_958_n953.n18 1.998
R12727 a_958_n953.n20 a_958_n953.n19 1.998
R12728 a_958_n953.n21 a_958_n953.n20 1.998
R12729 a_958_n953.n22 a_958_n953.n21 1.998
R12730 a_958_n953.n24 a_958_n953.n23 1.998
R12731 a_7272_n512.n0 a_7272_n512.t1 358.166
R12732 a_7272_n512.t4 a_7272_n512.t3 337.399
R12733 a_7272_n512.t3 a_7272_n512.t5 285.986
R12734 a_7272_n512.n0 a_7272_n512.t4 282.573
R12735 a_7272_n512.n1 a_7272_n512.t0 202.857
R12736 a_7272_n512.n1 a_7272_n512.n0 173.817
R12737 a_7272_n512.n1 a_7272_n512.t2 20.826
R12738 a_7272_n512.n2 a_7272_n512.n1 20.689
R12739 a_7177_n527.n0 a_7177_n527.t2 362.857
R12740 a_7177_n527.t3 a_7177_n527.t4 337.399
R12741 a_7177_n527.t4 a_7177_n527.t5 298.839
R12742 a_7177_n527.n0 a_7177_n527.t3 280.405
R12743 a_7177_n527.n1 a_7177_n527.t0 200
R12744 a_7177_n527.n1 a_7177_n527.n0 172.311
R12745 a_7177_n527.n2 a_7177_n527.n1 24
R12746 a_7177_n527.n1 a_7177_n527.t1 21.212
R12747 a_1317_4148.t0 a_1317_4148.t1 242.857
R12748 a_2577_2928.n0 a_2577_2928.t1 362.857
R12749 a_2577_2928.t3 a_2577_2928.t4 337.399
R12750 a_2577_2928.t4 a_2577_2928.t5 298.839
R12751 a_2577_2928.n0 a_2577_2928.t3 280.405
R12752 a_2577_2928.n1 a_2577_2928.t0 200
R12753 a_2577_2928.n1 a_2577_2928.n0 172.311
R12754 a_2577_2928.n2 a_2577_2928.n1 24
R12755 a_2577_2928.n1 a_2577_2928.t2 21.212
R12756 a_2672_2943.n0 a_2672_2943.t2 358.166
R12757 a_2672_2943.t5 a_2672_2943.t3 337.399
R12758 a_2672_2943.t3 a_2672_2943.t4 285.986
R12759 a_2672_2943.n0 a_2672_2943.t5 282.573
R12760 a_2672_2943.n1 a_2672_2943.t0 202.857
R12761 a_2672_2943.n1 a_2672_2943.n0 173.817
R12762 a_2672_2943.n1 a_2672_2943.t1 20.826
R12763 a_2672_2943.n2 a_2672_2943.n1 20.689
R12764 RWLB[6].n0 RWLB[6].t8 154.228
R12765 RWLB[6].n14 RWLB[6].t9 149.249
R12766 RWLB[6].n13 RWLB[6].t11 149.249
R12767 RWLB[6].n12 RWLB[6].t6 149.249
R12768 RWLB[6].n11 RWLB[6].t0 149.249
R12769 RWLB[6].n10 RWLB[6].t10 149.249
R12770 RWLB[6].n9 RWLB[6].t13 149.249
R12771 RWLB[6].n8 RWLB[6].t14 149.249
R12772 RWLB[6].n7 RWLB[6].t3 149.249
R12773 RWLB[6].n6 RWLB[6].t12 149.249
R12774 RWLB[6].n5 RWLB[6].t1 149.249
R12775 RWLB[6].n4 RWLB[6].t2 149.249
R12776 RWLB[6].n3 RWLB[6].t7 149.249
R12777 RWLB[6].n2 RWLB[6].t15 149.249
R12778 RWLB[6].n1 RWLB[6].t5 149.249
R12779 RWLB[6].n0 RWLB[6].t4 149.249
R12780 RWLB[6] RWLB[6].n14 47.816
R12781 RWLB[6].n1 RWLB[6].n0 4.979
R12782 RWLB[6].n2 RWLB[6].n1 4.979
R12783 RWLB[6].n3 RWLB[6].n2 4.979
R12784 RWLB[6].n4 RWLB[6].n3 4.979
R12785 RWLB[6].n5 RWLB[6].n4 4.979
R12786 RWLB[6].n6 RWLB[6].n5 4.979
R12787 RWLB[6].n7 RWLB[6].n6 4.979
R12788 RWLB[6].n8 RWLB[6].n7 4.979
R12789 RWLB[6].n9 RWLB[6].n8 4.979
R12790 RWLB[6].n10 RWLB[6].n9 4.979
R12791 RWLB[6].n11 RWLB[6].n10 4.979
R12792 RWLB[6].n12 RWLB[6].n11 4.979
R12793 RWLB[6].n13 RWLB[6].n12 4.979
R12794 RWLB[6].n14 RWLB[6].n13 4.979
R12795 a_2467_2180.t0 a_2467_2180.t1 242.857
R12796 a_2672_3666.n0 a_2672_3666.t1 358.166
R12797 a_2672_3666.t3 a_2672_3666.t4 337.399
R12798 a_2672_3666.t4 a_2672_3666.t5 285.986
R12799 a_2672_3666.n0 a_2672_3666.t3 282.573
R12800 a_2672_3666.n1 a_2672_3666.t0 202.857
R12801 a_2672_3666.n1 a_2672_3666.n0 173.817
R12802 a_2672_3666.n1 a_2672_3666.t2 20.826
R12803 a_2672_3666.n2 a_2672_3666.n1 20.689
R12804 a_2683_n953.n25 a_2683_n953.t27 561.971
R12805 a_2683_n953.n0 a_2683_n953.t21 461.908
R12806 a_2683_n953.t7 a_2683_n953.n25 108.635
R12807 a_2683_n953.n0 a_2683_n953.t22 79.512
R12808 a_2683_n953.n24 a_2683_n953.t26 65.401
R12809 a_2683_n953.n23 a_2683_n953.t10 65.401
R12810 a_2683_n953.n22 a_2683_n953.t2 65.401
R12811 a_2683_n953.n21 a_2683_n953.t19 65.401
R12812 a_2683_n953.n20 a_2683_n953.t14 65.401
R12813 a_2683_n953.n19 a_2683_n953.t9 65.401
R12814 a_2683_n953.n18 a_2683_n953.t24 65.401
R12815 a_2683_n953.n17 a_2683_n953.t5 65.401
R12816 a_2683_n953.n16 a_2683_n953.t23 65.401
R12817 a_2683_n953.n15 a_2683_n953.t3 65.401
R12818 a_2683_n953.n14 a_2683_n953.t12 65.401
R12819 a_2683_n953.n13 a_2683_n953.t0 65.401
R12820 a_2683_n953.n12 a_2683_n953.t8 65.401
R12821 a_2683_n953.n11 a_2683_n953.t16 65.401
R12822 a_2683_n953.n10 a_2683_n953.t6 65.401
R12823 a_2683_n953.n9 a_2683_n953.t13 65.401
R12824 a_2683_n953.n8 a_2683_n953.t11 65.401
R12825 a_2683_n953.n7 a_2683_n953.t25 65.401
R12826 a_2683_n953.n6 a_2683_n953.t1 65.401
R12827 a_2683_n953.n5 a_2683_n953.t17 65.401
R12828 a_2683_n953.n4 a_2683_n953.t4 65.401
R12829 a_2683_n953.n3 a_2683_n953.t15 65.401
R12830 a_2683_n953.n2 a_2683_n953.t18 65.401
R12831 a_2683_n953.n1 a_2683_n953.t20 65.401
R12832 a_2683_n953.n1 a_2683_n953.n0 5.64
R12833 a_2683_n953.n25 a_2683_n953.n24 4.438
R12834 a_2683_n953.n23 a_2683_n953.n22 2.524
R12835 a_2683_n953.n3 a_2683_n953.n2 2.498
R12836 a_2683_n953.n17 a_2683_n953.n16 2.364
R12837 a_2683_n953.n9 a_2683_n953.n8 2.355
R12838 a_2683_n953.n2 a_2683_n953.n1 1.998
R12839 a_2683_n953.n4 a_2683_n953.n3 1.998
R12840 a_2683_n953.n5 a_2683_n953.n4 1.998
R12841 a_2683_n953.n6 a_2683_n953.n5 1.998
R12842 a_2683_n953.n7 a_2683_n953.n6 1.998
R12843 a_2683_n953.n8 a_2683_n953.n7 1.998
R12844 a_2683_n953.n10 a_2683_n953.n9 1.998
R12845 a_2683_n953.n11 a_2683_n953.n10 1.998
R12846 a_2683_n953.n12 a_2683_n953.n11 1.998
R12847 a_2683_n953.n13 a_2683_n953.n12 1.998
R12848 a_2683_n953.n14 a_2683_n953.n13 1.998
R12849 a_2683_n953.n15 a_2683_n953.n14 1.998
R12850 a_2683_n953.n16 a_2683_n953.n15 1.998
R12851 a_2683_n953.n18 a_2683_n953.n17 1.998
R12852 a_2683_n953.n19 a_2683_n953.n18 1.998
R12853 a_2683_n953.n20 a_2683_n953.n19 1.998
R12854 a_2683_n953.n21 a_2683_n953.n20 1.998
R12855 a_2683_n953.n22 a_2683_n953.n21 1.998
R12856 a_2683_n953.n24 a_2683_n953.n23 1.998
R12857 a_7847_n271.n0 a_7847_n271.t2 358.166
R12858 a_7847_n271.t4 a_7847_n271.t5 337.399
R12859 a_7847_n271.t5 a_7847_n271.t3 285.986
R12860 a_7847_n271.n0 a_7847_n271.t4 282.573
R12861 a_7847_n271.n1 a_7847_n271.t0 202.857
R12862 a_7847_n271.n1 a_7847_n271.n0 173.817
R12863 a_7847_n271.n1 a_7847_n271.t1 20.826
R12864 a_7847_n271.n2 a_7847_n271.n1 20.689
R12865 a_8217_n271.t0 a_8217_n271.t1 242.857
R12866 a_7039_n8583.n0 a_7039_n8583.t4 1465.51
R12867 a_7039_n8583.n0 a_7039_n8583.t3 712.44
R12868 a_7039_n8583.n1 a_7039_n8583.t0 375.067
R12869 a_7039_n8583.n1 a_7039_n8583.t2 272.668
R12870 a_7039_n8583.n2 a_7039_n8583.n0 143.764
R12871 a_7039_n8583.t1 a_7039_n8583.n2 78.193
R12872 a_7039_n8583.n2 a_7039_n8583.n1 4.517
R12873 ADC9_OUT[3].n0 ADC9_OUT[3].t3 1355.37
R12874 ADC9_OUT[3].n0 ADC9_OUT[3].t4 820.859
R12875 ADC9_OUT[3].n3 ADC9_OUT[3].t0 326.879
R12876 ADC9_OUT[3].n2 ADC9_OUT[3].t2 266.644
R12877 ADC9_OUT[3].n1 ADC9_OUT[3].n0 149.035
R12878 ADC9_OUT[3].n3 ADC9_OUT[3].n2 57.223
R12879 ADC9_OUT[3].n1 ADC9_OUT[3].t1 45.968
R12880 ADC9_OUT[3] ADC9_OUT[3].n3 22.339
R12881 ADC9_OUT[3].n2 ADC9_OUT[3].n1 17.317
R12882 a_3266_n3770.n0 a_3266_n3770.t0 65.064
R12883 a_3266_n3770.n0 a_3266_n3770.t2 42.011
R12884 a_3266_n3770.t1 a_3266_n3770.n0 2.113
R12885 a_9008_n953.n25 a_9008_n953.t27 561.971
R12886 a_9008_n953.n0 a_9008_n953.t21 461.908
R12887 a_9008_n953.t6 a_9008_n953.n25 108.635
R12888 a_9008_n953.n0 a_9008_n953.t22 79.512
R12889 a_9008_n953.n24 a_9008_n953.t26 65.401
R12890 a_9008_n953.n23 a_9008_n953.t9 65.401
R12891 a_9008_n953.n22 a_9008_n953.t1 65.401
R12892 a_9008_n953.n21 a_9008_n953.t19 65.401
R12893 a_9008_n953.n20 a_9008_n953.t13 65.401
R12894 a_9008_n953.n19 a_9008_n953.t8 65.401
R12895 a_9008_n953.n18 a_9008_n953.t24 65.401
R12896 a_9008_n953.n17 a_9008_n953.t4 65.401
R12897 a_9008_n953.n16 a_9008_n953.t23 65.401
R12898 a_9008_n953.n15 a_9008_n953.t2 65.401
R12899 a_9008_n953.n14 a_9008_n953.t11 65.401
R12900 a_9008_n953.n13 a_9008_n953.t15 65.401
R12901 a_9008_n953.n12 a_9008_n953.t7 65.401
R12902 a_9008_n953.n11 a_9008_n953.t16 65.401
R12903 a_9008_n953.n10 a_9008_n953.t5 65.401
R12904 a_9008_n953.n9 a_9008_n953.t12 65.401
R12905 a_9008_n953.n8 a_9008_n953.t10 65.401
R12906 a_9008_n953.n7 a_9008_n953.t25 65.401
R12907 a_9008_n953.n6 a_9008_n953.t0 65.401
R12908 a_9008_n953.n5 a_9008_n953.t17 65.401
R12909 a_9008_n953.n4 a_9008_n953.t3 65.401
R12910 a_9008_n953.n3 a_9008_n953.t14 65.401
R12911 a_9008_n953.n2 a_9008_n953.t18 65.401
R12912 a_9008_n953.n1 a_9008_n953.t20 65.401
R12913 a_9008_n953.n1 a_9008_n953.n0 5.64
R12914 a_9008_n953.n25 a_9008_n953.n24 4.438
R12915 a_9008_n953.n23 a_9008_n953.n22 2.524
R12916 a_9008_n953.n3 a_9008_n953.n2 2.498
R12917 a_9008_n953.n17 a_9008_n953.n16 2.364
R12918 a_9008_n953.n9 a_9008_n953.n8 2.355
R12919 a_9008_n953.n2 a_9008_n953.n1 1.998
R12920 a_9008_n953.n4 a_9008_n953.n3 1.998
R12921 a_9008_n953.n5 a_9008_n953.n4 1.998
R12922 a_9008_n953.n6 a_9008_n953.n5 1.998
R12923 a_9008_n953.n7 a_9008_n953.n6 1.998
R12924 a_9008_n953.n8 a_9008_n953.n7 1.998
R12925 a_9008_n953.n10 a_9008_n953.n9 1.998
R12926 a_9008_n953.n11 a_9008_n953.n10 1.998
R12927 a_9008_n953.n12 a_9008_n953.n11 1.998
R12928 a_9008_n953.n13 a_9008_n953.n12 1.998
R12929 a_9008_n953.n14 a_9008_n953.n13 1.998
R12930 a_9008_n953.n15 a_9008_n953.n14 1.998
R12931 a_9008_n953.n16 a_9008_n953.n15 1.998
R12932 a_9008_n953.n18 a_9008_n953.n17 1.998
R12933 a_9008_n953.n19 a_9008_n953.n18 1.998
R12934 a_9008_n953.n20 a_9008_n953.n19 1.998
R12935 a_9008_n953.n21 a_9008_n953.n20 1.998
R12936 a_9008_n953.n22 a_9008_n953.n21 1.998
R12937 a_9008_n953.n24 a_9008_n953.n23 1.998
R12938 a_9078_n2086.t0 a_9078_n2086.t1 34.8
R12939 a_8422_n812.n0 a_8422_n812.t1 358.166
R12940 a_8422_n812.t5 a_8422_n812.t4 337.399
R12941 a_8422_n812.t4 a_8422_n812.t3 285.986
R12942 a_8422_n812.n0 a_8422_n812.t5 282.573
R12943 a_8422_n812.n1 a_8422_n812.t0 202.857
R12944 a_8422_n812.n1 a_8422_n812.n0 173.817
R12945 a_8422_n812.n1 a_8422_n812.t2 20.826
R12946 a_8422_n812.n2 a_8422_n812.n1 20.689
R12947 a_8792_n812.t0 a_8792_n812.t1 242.857
R12948 a_4972_1457.n0 a_4972_1457.t1 358.166
R12949 a_4972_1457.t3 a_4972_1457.t5 337.399
R12950 a_4972_1457.t5 a_4972_1457.t4 285.986
R12951 a_4972_1457.n0 a_4972_1457.t3 282.573
R12952 a_4972_1457.n1 a_4972_1457.t0 202.857
R12953 a_4972_1457.n1 a_4972_1457.n0 173.817
R12954 a_4972_1457.n1 a_4972_1457.t2 20.826
R12955 a_4972_1457.n2 a_4972_1457.n1 20.689
R12956 a_4877_1442.n0 a_4877_1442.t2 362.857
R12957 a_4877_1442.t4 a_4877_1442.t3 337.399
R12958 a_4877_1442.t3 a_4877_1442.t5 298.839
R12959 a_4877_1442.n0 a_4877_1442.t4 280.405
R12960 a_4877_1442.n1 a_4877_1442.t0 200
R12961 a_4877_1442.n1 a_4877_1442.n0 172.311
R12962 a_4877_1442.n2 a_4877_1442.n1 24
R12963 a_4877_1442.n1 a_4877_1442.t1 21.212
R12964 a_3727_n45.n0 a_3727_n45.t2 362.857
R12965 a_3727_n45.t4 a_3727_n45.t3 337.399
R12966 a_3727_n45.t3 a_3727_n45.t5 298.839
R12967 a_3727_n45.n0 a_3727_n45.t4 280.405
R12968 a_3727_n45.n1 a_3727_n45.t0 200
R12969 a_3727_n45.n1 a_3727_n45.n0 172.311
R12970 a_3727_n45.n2 a_3727_n45.n1 24
R12971 a_3727_n45.n1 a_3727_n45.t1 21.212
R12972 a_3822_n30.n0 a_3822_n30.t2 358.166
R12973 a_3822_n30.t3 a_3822_n30.t5 337.399
R12974 a_3822_n30.t5 a_3822_n30.t4 285.986
R12975 a_3822_n30.n0 a_3822_n30.t3 282.573
R12976 a_3822_n30.n1 a_3822_n30.t0 202.857
R12977 a_3822_n30.n1 a_3822_n30.n0 173.817
R12978 a_3822_n30.n1 a_3822_n30.t1 20.826
R12979 a_3822_n30.n2 a_3822_n30.n1 20.689
R12980 Iref1.n0 Iref1.t7 464.674
R12981 Iref1.n14 Iref1.t6 457.028
R12982 Iref1.n13 Iref1.t15 457.028
R12983 Iref1.n12 Iref1.t8 457.028
R12984 Iref1.n10 Iref1.t13 457.028
R12985 Iref1.n9 Iref1.t1 457.028
R12986 Iref1.n8 Iref1.t4 457.028
R12987 Iref1.n7 Iref1.t11 457.028
R12988 Iref1.n6 Iref1.t3 457.028
R12989 Iref1.n5 Iref1.t10 457.028
R12990 Iref1.n4 Iref1.t2 457.028
R12991 Iref1.n3 Iref1.t9 457.028
R12992 Iref1.n2 Iref1.t12 457.028
R12993 Iref1.n0 Iref1.t0 457.028
R12994 Iref1.n11 Iref1.t14 456.275
R12995 Iref1.n1 Iref1.t5 454.769
R12996 Iref1 Iref1.n14 39.35
R12997 Iref1.n12 Iref1.n11 8.671
R12998 Iref1.n13 Iref1.n12 8.671
R12999 Iref1.n10 Iref1.n9 8.649
R13000 Iref1.n11 Iref1.n10 8.649
R13001 Iref1.n1 Iref1.n0 8.634
R13002 Iref1.n4 Iref1.n3 8.634
R13003 Iref1.n5 Iref1.n4 8.634
R13004 Iref1.n6 Iref1.n5 8.634
R13005 Iref1.n7 Iref1.n6 8.634
R13006 Iref1.n8 Iref1.n7 8.634
R13007 Iref1.n9 Iref1.n8 8.634
R13008 Iref1.n2 Iref1.n1 8.627
R13009 Iref1.n3 Iref1.n2 8.627
R13010 Iref1.n14 Iref1.n13 6.568
R13011 a_n2148_n5293.t1 a_n2148_n5293.t0 336.814
R13012 a_n2207_n5338.t0 a_n2207_n5338.t1 68.74
R13013 a_372_3666.n0 a_372_3666.t2 358.166
R13014 a_372_3666.t4 a_372_3666.t3 337.399
R13015 a_372_3666.t3 a_372_3666.t5 285.986
R13016 a_372_3666.n0 a_372_3666.t4 282.573
R13017 a_372_3666.n1 a_372_3666.t0 202.857
R13018 a_372_3666.n1 a_372_3666.n0 173.817
R13019 a_372_3666.n1 a_372_3666.t1 20.826
R13020 a_372_3666.n2 a_372_3666.n1 20.689
R13021 a_277_3651.n0 a_277_3651.t1 362.857
R13022 a_277_3651.t5 a_277_3651.t3 337.399
R13023 a_277_3651.t3 a_277_3651.t4 298.839
R13024 a_277_3651.n0 a_277_3651.t5 280.405
R13025 a_277_3651.n1 a_277_3651.t2 200
R13026 a_277_3651.n1 a_277_3651.n0 172.311
R13027 a_277_3651.n2 a_277_3651.n1 24
R13028 a_277_3651.n1 a_277_3651.t0 21.212
R13029 a_1427_n1068.n0 a_1427_n1068.t0 362.857
R13030 a_1427_n1068.t3 a_1427_n1068.t4 337.399
R13031 a_1427_n1068.t4 a_1427_n1068.t5 298.839
R13032 a_1427_n1068.n0 a_1427_n1068.t3 280.405
R13033 a_1427_n1068.n1 a_1427_n1068.t1 200
R13034 a_1427_n1068.n1 a_1427_n1068.n0 172.311
R13035 a_1427_n1068.n2 a_1427_n1068.n1 24
R13036 a_1427_n1068.n1 a_1427_n1068.t2 21.212
R13037 a_1522_n1053.n0 a_1522_n1053.t1 358.166
R13038 a_1522_n1053.t4 a_1522_n1053.t3 337.399
R13039 a_1522_n1053.t3 a_1522_n1053.t5 285.986
R13040 a_1522_n1053.n0 a_1522_n1053.t4 282.573
R13041 a_1522_n1053.n1 a_1522_n1053.t2 202.857
R13042 a_1522_n1053.n1 a_1522_n1053.n0 173.817
R13043 a_1522_n1053.n1 a_1522_n1053.t0 20.826
R13044 a_1522_n1053.n2 a_1522_n1053.n1 20.689
R13045 a_13033_n7203.n0 a_13033_n7203.t0 63.08
R13046 a_13033_n7203.n0 a_13033_n7203.t2 41.305
R13047 a_13033_n7203.t1 a_13033_n7203.n0 2.251
R13048 a_13171_n7203.t1 a_13171_n7203.t0 68.741
R13049 a_6602_2647.n0 a_6602_2647.t1 362.857
R13050 a_6602_2647.t4 a_6602_2647.t3 337.399
R13051 a_6602_2647.t3 a_6602_2647.t5 298.839
R13052 a_6602_2647.n0 a_6602_2647.t4 280.405
R13053 a_6602_2647.n1 a_6602_2647.t0 200
R13054 a_6602_2647.n1 a_6602_2647.n0 172.311
R13055 a_6602_2647.n2 a_6602_2647.n1 24
R13056 a_6602_2647.n1 a_6602_2647.t2 21.212
R13057 a_6697_2662.n0 a_6697_2662.t1 358.166
R13058 a_6697_2662.t3 a_6697_2662.t4 337.399
R13059 a_6697_2662.t4 a_6697_2662.t5 285.986
R13060 a_6697_2662.n0 a_6697_2662.t3 282.573
R13061 a_6697_2662.n1 a_6697_2662.t2 202.857
R13062 a_6697_2662.n1 a_6697_2662.n0 173.817
R13063 a_6697_2662.n1 a_6697_2662.t0 20.826
R13064 a_6697_2662.n2 a_6697_2662.n1 20.689
R13065 a_8997_1457.n0 a_8997_1457.t1 358.166
R13066 a_8997_1457.t4 a_8997_1457.t5 337.399
R13067 a_8997_1457.t5 a_8997_1457.t3 285.986
R13068 a_8997_1457.n0 a_8997_1457.t4 282.573
R13069 a_8997_1457.n1 a_8997_1457.t2 202.857
R13070 a_8997_1457.n1 a_8997_1457.n0 173.817
R13071 a_8997_1457.n1 a_8997_1457.t0 20.826
R13072 a_8997_1457.n2 a_8997_1457.n1 20.689
R13073 a_9367_1457.t0 a_9367_1457.t1 242.857
R13074 WWLD[4].n0 WWLD[4].t14 262.032
R13075 WWLD[4].n29 WWLD[4].t17 260.715
R13076 WWLD[4].n27 WWLD[4].t19 260.715
R13077 WWLD[4].n25 WWLD[4].t7 260.715
R13078 WWLD[4].n23 WWLD[4].t30 260.715
R13079 WWLD[4].n21 WWLD[4].t9 260.715
R13080 WWLD[4].n19 WWLD[4].t25 260.715
R13081 WWLD[4].n17 WWLD[4].t16 260.715
R13082 WWLD[4].n15 WWLD[4].t3 260.715
R13083 WWLD[4].n13 WWLD[4].t21 260.715
R13084 WWLD[4].n11 WWLD[4].t31 260.715
R13085 WWLD[4].n9 WWLD[4].t18 260.715
R13086 WWLD[4].n7 WWLD[4].t5 260.715
R13087 WWLD[4].n5 WWLD[4].t26 260.715
R13088 WWLD[4].n3 WWLD[4].t10 260.715
R13089 WWLD[4].n1 WWLD[4].t22 260.715
R13090 WWLD[4].n30 WWLD[4].t20 259.254
R13091 WWLD[4].n28 WWLD[4].t29 259.254
R13092 WWLD[4].n26 WWLD[4].t8 259.254
R13093 WWLD[4].n24 WWLD[4].t23 259.254
R13094 WWLD[4].n22 WWLD[4].t13 259.254
R13095 WWLD[4].n20 WWLD[4].t0 259.254
R13096 WWLD[4].n18 WWLD[4].t11 259.254
R13097 WWLD[4].n16 WWLD[4].t27 259.254
R13098 WWLD[4].n14 WWLD[4].t15 259.254
R13099 WWLD[4].n12 WWLD[4].t4 259.254
R13100 WWLD[4].n10 WWLD[4].t24 259.254
R13101 WWLD[4].n8 WWLD[4].t1 259.254
R13102 WWLD[4].n6 WWLD[4].t2 259.254
R13103 WWLD[4].n4 WWLD[4].t6 259.254
R13104 WWLD[4].n2 WWLD[4].t28 259.254
R13105 WWLD[4].n0 WWLD[4].t12 259.254
R13106 WWLD[4] WWLD[4].n30 44.647
R13107 WWLD[4].n1 WWLD[4].n0 3.576
R13108 WWLD[4].n3 WWLD[4].n2 3.576
R13109 WWLD[4].n5 WWLD[4].n4 3.576
R13110 WWLD[4].n7 WWLD[4].n6 3.576
R13111 WWLD[4].n9 WWLD[4].n8 3.576
R13112 WWLD[4].n11 WWLD[4].n10 3.576
R13113 WWLD[4].n13 WWLD[4].n12 3.576
R13114 WWLD[4].n15 WWLD[4].n14 3.576
R13115 WWLD[4].n17 WWLD[4].n16 3.576
R13116 WWLD[4].n19 WWLD[4].n18 3.576
R13117 WWLD[4].n21 WWLD[4].n20 3.576
R13118 WWLD[4].n23 WWLD[4].n22 3.576
R13119 WWLD[4].n25 WWLD[4].n24 3.576
R13120 WWLD[4].n27 WWLD[4].n26 3.576
R13121 WWLD[4].n29 WWLD[4].n28 3.576
R13122 WWLD[4].n2 WWLD[4].n1 1.317
R13123 WWLD[4].n4 WWLD[4].n3 1.317
R13124 WWLD[4].n6 WWLD[4].n5 1.317
R13125 WWLD[4].n8 WWLD[4].n7 1.317
R13126 WWLD[4].n10 WWLD[4].n9 1.317
R13127 WWLD[4].n12 WWLD[4].n11 1.317
R13128 WWLD[4].n14 WWLD[4].n13 1.317
R13129 WWLD[4].n16 WWLD[4].n15 1.317
R13130 WWLD[4].n18 WWLD[4].n17 1.317
R13131 WWLD[4].n20 WWLD[4].n19 1.317
R13132 WWLD[4].n22 WWLD[4].n21 1.317
R13133 WWLD[4].n24 WWLD[4].n23 1.317
R13134 WWLD[4].n26 WWLD[4].n25 1.317
R13135 WWLD[4].n28 WWLD[4].n27 1.317
R13136 WWLD[4].n30 WWLD[4].n29 1.317
R13137 a_3247_n271.n0 a_3247_n271.t1 358.166
R13138 a_3247_n271.t4 a_3247_n271.t5 337.399
R13139 a_3247_n271.t5 a_3247_n271.t3 285.986
R13140 a_3247_n271.n0 a_3247_n271.t4 282.573
R13141 a_3247_n271.n1 a_3247_n271.t0 202.857
R13142 a_3247_n271.n1 a_3247_n271.n0 173.817
R13143 a_3247_n271.n1 a_3247_n271.t2 20.826
R13144 a_3247_n271.n2 a_3247_n271.n1 20.689
R13145 a_8902_n827.n0 a_8902_n827.t1 362.857
R13146 a_8902_n827.t3 a_8902_n827.t5 337.399
R13147 a_8902_n827.t5 a_8902_n827.t4 298.839
R13148 a_8902_n827.n0 a_8902_n827.t3 280.405
R13149 a_8902_n827.n1 a_8902_n827.t0 200
R13150 a_8902_n827.n1 a_8902_n827.n0 172.311
R13151 a_8902_n827.n2 a_8902_n827.n1 24
R13152 a_8902_n827.n1 a_8902_n827.t2 21.212
R13153 a_8997_n812.n0 a_8997_n812.t1 358.166
R13154 a_8997_n812.t4 a_8997_n812.t5 337.399
R13155 a_8997_n812.t5 a_8997_n812.t3 285.986
R13156 a_8997_n812.n0 a_8997_n812.t4 282.573
R13157 a_8997_n812.n1 a_8997_n812.t2 202.857
R13158 a_8997_n812.n1 a_8997_n812.n0 173.817
R13159 a_8997_n812.n1 a_8997_n812.t0 20.826
R13160 a_8997_n812.n2 a_8997_n812.n1 20.689
R13161 WWLD[1].n0 WWLD[1].t15 262.032
R13162 WWLD[1].n29 WWLD[1].t18 260.715
R13163 WWLD[1].n27 WWLD[1].t21 260.715
R13164 WWLD[1].n25 WWLD[1].t3 260.715
R13165 WWLD[1].n23 WWLD[1].t29 260.715
R13166 WWLD[1].n21 WWLD[1].t9 260.715
R13167 WWLD[1].n19 WWLD[1].t26 260.715
R13168 WWLD[1].n17 WWLD[1].t17 260.715
R13169 WWLD[1].n15 WWLD[1].t0 260.715
R13170 WWLD[1].n13 WWLD[1].t22 260.715
R13171 WWLD[1].n11 WWLD[1].t30 260.715
R13172 WWLD[1].n9 WWLD[1].t19 260.715
R13173 WWLD[1].n7 WWLD[1].t1 260.715
R13174 WWLD[1].n5 WWLD[1].t27 260.715
R13175 WWLD[1].n3 WWLD[1].t10 260.715
R13176 WWLD[1].n1 WWLD[1].t23 260.715
R13177 WWLD[1].n30 WWLD[1].t2 259.254
R13178 WWLD[1].n28 WWLD[1].t8 259.254
R13179 WWLD[1].n26 WWLD[1].t20 259.254
R13180 WWLD[1].n24 WWLD[1].t4 259.254
R13181 WWLD[1].n22 WWLD[1].t28 259.254
R13182 WWLD[1].n20 WWLD[1].t11 259.254
R13183 WWLD[1].n18 WWLD[1].t24 259.254
R13184 WWLD[1].n16 WWLD[1].t6 259.254
R13185 WWLD[1].n14 WWLD[1].t31 259.254
R13186 WWLD[1].n12 WWLD[1].t14 259.254
R13187 WWLD[1].n10 WWLD[1].t5 259.254
R13188 WWLD[1].n8 WWLD[1].t12 259.254
R13189 WWLD[1].n6 WWLD[1].t13 259.254
R13190 WWLD[1].n4 WWLD[1].t16 259.254
R13191 WWLD[1].n2 WWLD[1].t7 259.254
R13192 WWLD[1].n0 WWLD[1].t25 259.254
R13193 WWLD[1] WWLD[1].n30 44.647
R13194 WWLD[1].n1 WWLD[1].n0 3.576
R13195 WWLD[1].n3 WWLD[1].n2 3.576
R13196 WWLD[1].n5 WWLD[1].n4 3.576
R13197 WWLD[1].n7 WWLD[1].n6 3.576
R13198 WWLD[1].n9 WWLD[1].n8 3.576
R13199 WWLD[1].n11 WWLD[1].n10 3.576
R13200 WWLD[1].n13 WWLD[1].n12 3.576
R13201 WWLD[1].n15 WWLD[1].n14 3.576
R13202 WWLD[1].n17 WWLD[1].n16 3.576
R13203 WWLD[1].n19 WWLD[1].n18 3.576
R13204 WWLD[1].n21 WWLD[1].n20 3.576
R13205 WWLD[1].n23 WWLD[1].n22 3.576
R13206 WWLD[1].n25 WWLD[1].n24 3.576
R13207 WWLD[1].n27 WWLD[1].n26 3.576
R13208 WWLD[1].n29 WWLD[1].n28 3.576
R13209 WWLD[1].n2 WWLD[1].n1 1.317
R13210 WWLD[1].n4 WWLD[1].n3 1.317
R13211 WWLD[1].n6 WWLD[1].n5 1.317
R13212 WWLD[1].n8 WWLD[1].n7 1.317
R13213 WWLD[1].n10 WWLD[1].n9 1.317
R13214 WWLD[1].n12 WWLD[1].n11 1.317
R13215 WWLD[1].n14 WWLD[1].n13 1.317
R13216 WWLD[1].n16 WWLD[1].n15 1.317
R13217 WWLD[1].n18 WWLD[1].n17 1.317
R13218 WWLD[1].n20 WWLD[1].n19 1.317
R13219 WWLD[1].n22 WWLD[1].n21 1.317
R13220 WWLD[1].n24 WWLD[1].n23 1.317
R13221 WWLD[1].n26 WWLD[1].n25 1.317
R13222 WWLD[1].n28 WWLD[1].n27 1.317
R13223 WWLD[1].n30 WWLD[1].n29 1.317
R13224 a_4302_4430.n0 a_4302_4430.t1 362.857
R13225 a_4302_4430.t3 a_4302_4430.t5 337.399
R13226 a_4302_4430.t5 a_4302_4430.t4 298.839
R13227 a_4302_4430.n0 a_4302_4430.t3 280.405
R13228 a_4302_4430.n1 a_4302_4430.t0 200
R13229 a_4302_4430.n1 a_4302_4430.n0 172.311
R13230 a_4302_4430.n2 a_4302_4430.n1 24
R13231 a_4302_4430.n1 a_4302_4430.t2 21.212
R13232 a_7847_3425.n0 a_7847_3425.t2 358.166
R13233 a_7847_3425.t4 a_7847_3425.t5 337.399
R13234 a_7847_3425.t5 a_7847_3425.t3 285.986
R13235 a_7847_3425.n0 a_7847_3425.t4 282.573
R13236 a_7847_3425.n1 a_7847_3425.t0 202.857
R13237 a_7847_3425.n1 a_7847_3425.n0 173.817
R13238 a_7847_3425.n1 a_7847_3425.t1 20.826
R13239 a_7847_3425.n2 a_7847_3425.n1 20.689
R13240 a_8217_3425.t0 a_8217_3425.t1 242.857
R13241 a_6697_3907.n0 a_6697_3907.t1 358.166
R13242 a_6697_3907.t4 a_6697_3907.t5 337.399
R13243 a_6697_3907.t5 a_6697_3907.t3 285.986
R13244 a_6697_3907.n0 a_6697_3907.t4 282.573
R13245 a_6697_3907.n1 a_6697_3907.t2 202.857
R13246 a_6697_3907.n1 a_6697_3907.n0 173.817
R13247 a_6697_3907.n1 a_6697_3907.t0 20.826
R13248 a_6697_3907.n2 a_6697_3907.n1 20.689
R13249 a_6708_n953.n25 a_6708_n953.t27 561.971
R13250 a_6708_n953.n0 a_6708_n953.t22 461.908
R13251 a_6708_n953.t6 a_6708_n953.n25 108.635
R13252 a_6708_n953.n0 a_6708_n953.t23 79.512
R13253 a_6708_n953.n24 a_6708_n953.t24 65.401
R13254 a_6708_n953.n23 a_6708_n953.t10 65.401
R13255 a_6708_n953.n22 a_6708_n953.t2 65.401
R13256 a_6708_n953.n21 a_6708_n953.t7 65.401
R13257 a_6708_n953.n20 a_6708_n953.t14 65.401
R13258 a_6708_n953.n19 a_6708_n953.t9 65.401
R13259 a_6708_n953.n18 a_6708_n953.t21 65.401
R13260 a_6708_n953.n17 a_6708_n953.t5 65.401
R13261 a_6708_n953.n16 a_6708_n953.t26 65.401
R13262 a_6708_n953.n15 a_6708_n953.t3 65.401
R13263 a_6708_n953.n14 a_6708_n953.t12 65.401
R13264 a_6708_n953.n13 a_6708_n953.t15 65.401
R13265 a_6708_n953.n12 a_6708_n953.t8 65.401
R13266 a_6708_n953.n11 a_6708_n953.t18 65.401
R13267 a_6708_n953.n10 a_6708_n953.t1 65.401
R13268 a_6708_n953.n9 a_6708_n953.t13 65.401
R13269 a_6708_n953.n8 a_6708_n953.t11 65.401
R13270 a_6708_n953.n7 a_6708_n953.t25 65.401
R13271 a_6708_n953.n6 a_6708_n953.t0 65.401
R13272 a_6708_n953.n5 a_6708_n953.t19 65.401
R13273 a_6708_n953.n4 a_6708_n953.t4 65.401
R13274 a_6708_n953.n3 a_6708_n953.t16 65.401
R13275 a_6708_n953.n2 a_6708_n953.t17 65.401
R13276 a_6708_n953.n1 a_6708_n953.t20 65.401
R13277 a_6708_n953.n1 a_6708_n953.n0 5.64
R13278 a_6708_n953.n25 a_6708_n953.n24 4.438
R13279 a_6708_n953.n23 a_6708_n953.n22 2.524
R13280 a_6708_n953.n3 a_6708_n953.n2 2.498
R13281 a_6708_n953.n17 a_6708_n953.n16 2.364
R13282 a_6708_n953.n9 a_6708_n953.n8 2.355
R13283 a_6708_n953.n2 a_6708_n953.n1 1.998
R13284 a_6708_n953.n4 a_6708_n953.n3 1.998
R13285 a_6708_n953.n5 a_6708_n953.n4 1.998
R13286 a_6708_n953.n6 a_6708_n953.n5 1.998
R13287 a_6708_n953.n7 a_6708_n953.n6 1.998
R13288 a_6708_n953.n8 a_6708_n953.n7 1.998
R13289 a_6708_n953.n10 a_6708_n953.n9 1.998
R13290 a_6708_n953.n11 a_6708_n953.n10 1.998
R13291 a_6708_n953.n12 a_6708_n953.n11 1.998
R13292 a_6708_n953.n13 a_6708_n953.n12 1.998
R13293 a_6708_n953.n14 a_6708_n953.n13 1.998
R13294 a_6708_n953.n15 a_6708_n953.n14 1.998
R13295 a_6708_n953.n16 a_6708_n953.n15 1.998
R13296 a_6708_n953.n18 a_6708_n953.n17 1.998
R13297 a_6708_n953.n19 a_6708_n953.n18 1.998
R13298 a_6708_n953.n20 a_6708_n953.n19 1.998
R13299 a_6708_n953.n21 a_6708_n953.n20 1.998
R13300 a_6708_n953.n22 a_6708_n953.n21 1.998
R13301 a_6708_n953.n24 a_6708_n953.n23 1.998
R13302 RWLB[11].n0 RWLB[11].t5 154.228
R13303 RWLB[11].n14 RWLB[11].t10 149.249
R13304 RWLB[11].n13 RWLB[11].t9 149.249
R13305 RWLB[11].n12 RWLB[11].t1 149.249
R13306 RWLB[11].n11 RWLB[11].t13 149.249
R13307 RWLB[11].n10 RWLB[11].t4 149.249
R13308 RWLB[11].n9 RWLB[11].t3 149.249
R13309 RWLB[11].n8 RWLB[11].t7 149.249
R13310 RWLB[11].n7 RWLB[11].t6 149.249
R13311 RWLB[11].n6 RWLB[11].t15 149.249
R13312 RWLB[11].n5 RWLB[11].t14 149.249
R13313 RWLB[11].n4 RWLB[11].t0 149.249
R13314 RWLB[11].n3 RWLB[11].t11 149.249
R13315 RWLB[11].n2 RWLB[11].t8 149.249
R13316 RWLB[11].n1 RWLB[11].t2 149.249
R13317 RWLB[11].n0 RWLB[11].t12 149.249
R13318 RWLB[11] RWLB[11].n14 47.816
R13319 RWLB[11].n1 RWLB[11].n0 4.979
R13320 RWLB[11].n2 RWLB[11].n1 4.979
R13321 RWLB[11].n3 RWLB[11].n2 4.979
R13322 RWLB[11].n4 RWLB[11].n3 4.979
R13323 RWLB[11].n5 RWLB[11].n4 4.979
R13324 RWLB[11].n6 RWLB[11].n5 4.979
R13325 RWLB[11].n7 RWLB[11].n6 4.979
R13326 RWLB[11].n8 RWLB[11].n7 4.979
R13327 RWLB[11].n9 RWLB[11].n8 4.979
R13328 RWLB[11].n10 RWLB[11].n9 4.979
R13329 RWLB[11].n11 RWLB[11].n10 4.979
R13330 RWLB[11].n12 RWLB[11].n11 4.979
R13331 RWLB[11].n13 RWLB[11].n12 4.979
R13332 RWLB[11].n14 RWLB[11].n13 4.979
R13333 a_6040_n953.t36 a_6040_n953.n46 176.385
R13334 a_6040_n953.n22 a_6040_n953.t11 67.378
R13335 a_6040_n953.n0 a_6040_n953.t15 66.92
R13336 a_6040_n953.n1 a_6040_n953.t13 66.92
R13337 a_6040_n953.n2 a_6040_n953.t4 66.92
R13338 a_6040_n953.n3 a_6040_n953.t12 66.92
R13339 a_6040_n953.n4 a_6040_n953.t0 66.92
R13340 a_6040_n953.n5 a_6040_n953.t48 66.92
R13341 a_6040_n953.n6 a_6040_n953.t42 66.92
R13342 a_6040_n953.n7 a_6040_n953.t46 66.92
R13343 a_6040_n953.n8 a_6040_n953.t24 66.92
R13344 a_6040_n953.n9 a_6040_n953.t30 66.92
R13345 a_6040_n953.n10 a_6040_n953.t18 66.92
R13346 a_6040_n953.n11 a_6040_n953.t33 66.92
R13347 a_6040_n953.n12 a_6040_n953.t28 66.92
R13348 a_6040_n953.n13 a_6040_n953.t44 66.92
R13349 a_6040_n953.n14 a_6040_n953.t47 66.92
R13350 a_6040_n953.n15 a_6040_n953.t45 66.92
R13351 a_6040_n953.n16 a_6040_n953.t17 66.92
R13352 a_6040_n953.n17 a_6040_n953.t26 66.92
R13353 a_6040_n953.n18 a_6040_n953.t21 66.92
R13354 a_6040_n953.n19 a_6040_n953.t27 66.92
R13355 a_6040_n953.n20 a_6040_n953.t8 66.92
R13356 a_6040_n953.n21 a_6040_n953.t3 66.92
R13357 a_6040_n953.n22 a_6040_n953.t6 66.92
R13358 a_6040_n953.n23 a_6040_n953.t1 65.518
R13359 a_6040_n953.n45 a_6040_n953.t14 63.519
R13360 a_6040_n953.n44 a_6040_n953.t10 63.519
R13361 a_6040_n953.n43 a_6040_n953.t16 63.519
R13362 a_6040_n953.n42 a_6040_n953.t2 63.519
R13363 a_6040_n953.n41 a_6040_n953.t37 63.519
R13364 a_6040_n953.n40 a_6040_n953.t41 63.519
R13365 a_6040_n953.n39 a_6040_n953.t20 63.519
R13366 a_6040_n953.n38 a_6040_n953.t19 63.519
R13367 a_6040_n953.n37 a_6040_n953.t22 63.519
R13368 a_6040_n953.n36 a_6040_n953.t40 63.519
R13369 a_6040_n953.n35 a_6040_n953.t32 63.519
R13370 a_6040_n953.n34 a_6040_n953.t34 63.519
R13371 a_6040_n953.n33 a_6040_n953.t38 63.519
R13372 a_6040_n953.n32 a_6040_n953.t23 63.519
R13373 a_6040_n953.n31 a_6040_n953.t43 63.519
R13374 a_6040_n953.n30 a_6040_n953.t39 63.519
R13375 a_6040_n953.n29 a_6040_n953.t35 63.519
R13376 a_6040_n953.n28 a_6040_n953.t31 63.519
R13377 a_6040_n953.n27 a_6040_n953.t29 63.519
R13378 a_6040_n953.n26 a_6040_n953.t25 63.519
R13379 a_6040_n953.n25 a_6040_n953.t7 63.519
R13380 a_6040_n953.n24 a_6040_n953.t9 63.519
R13381 a_6040_n953.n23 a_6040_n953.t5 63.519
R13382 a_6040_n953.n46 a_6040_n953.n0 19.599
R13383 a_6040_n953.n46 a_6040_n953.n45 15.67
R13384 a_6040_n953.n44 a_6040_n953.n43 2.524
R13385 a_6040_n953.n24 a_6040_n953.n23 2.498
R13386 a_6040_n953.n21 a_6040_n953.n22 2.495
R13387 a_6040_n953.n1 a_6040_n953.n2 2.459
R13388 a_6040_n953.n38 a_6040_n953.n37 2.364
R13389 a_6040_n953.n30 a_6040_n953.n29 2.355
R13390 a_6040_n953.n7 a_6040_n953.n8 2.299
R13391 a_6040_n953.n15 a_6040_n953.n16 2.29
R13392 a_6040_n953.n16 a_6040_n953.n17 2.057
R13393 a_6040_n953.n8 a_6040_n953.n9 2.057
R13394 a_6040_n953.n2 a_6040_n953.n3 2.057
R13395 a_6040_n953.n0 a_6040_n953.n1 2.057
R13396 a_6040_n953.n45 a_6040_n953.n44 1.998
R13397 a_6040_n953.n43 a_6040_n953.n42 1.998
R13398 a_6040_n953.n42 a_6040_n953.n41 1.998
R13399 a_6040_n953.n41 a_6040_n953.n40 1.998
R13400 a_6040_n953.n40 a_6040_n953.n39 1.998
R13401 a_6040_n953.n39 a_6040_n953.n38 1.998
R13402 a_6040_n953.n37 a_6040_n953.n36 1.998
R13403 a_6040_n953.n36 a_6040_n953.n35 1.998
R13404 a_6040_n953.n35 a_6040_n953.n34 1.998
R13405 a_6040_n953.n34 a_6040_n953.n33 1.998
R13406 a_6040_n953.n33 a_6040_n953.n32 1.998
R13407 a_6040_n953.n32 a_6040_n953.n31 1.998
R13408 a_6040_n953.n31 a_6040_n953.n30 1.998
R13409 a_6040_n953.n29 a_6040_n953.n28 1.998
R13410 a_6040_n953.n28 a_6040_n953.n27 1.998
R13411 a_6040_n953.n27 a_6040_n953.n26 1.998
R13412 a_6040_n953.n26 a_6040_n953.n25 1.998
R13413 a_6040_n953.n25 a_6040_n953.n24 1.998
R13414 a_6040_n953.n20 a_6040_n953.n21 1.995
R13415 a_6040_n953.n19 a_6040_n953.n20 1.995
R13416 a_6040_n953.n18 a_6040_n953.n19 1.995
R13417 a_6040_n953.n17 a_6040_n953.n18 1.995
R13418 a_6040_n953.n14 a_6040_n953.n15 1.995
R13419 a_6040_n953.n13 a_6040_n953.n14 1.995
R13420 a_6040_n953.n12 a_6040_n953.n13 1.995
R13421 a_6040_n953.n11 a_6040_n953.n12 1.995
R13422 a_6040_n953.n10 a_6040_n953.n11 1.995
R13423 a_6040_n953.n9 a_6040_n953.n10 1.995
R13424 a_6040_n953.n6 a_6040_n953.n7 1.995
R13425 a_6040_n953.n5 a_6040_n953.n6 1.995
R13426 a_6040_n953.n4 a_6040_n953.n5 1.995
R13427 a_6040_n953.n3 a_6040_n953.n4 1.995
R13428 a_6492_975.t0 a_6492_975.t1 242.857
R13429 a_8340_4445.t0 a_8340_4445.t1 242.857
R13430 WWL[11].n0 WWL[11].t14 262.032
R13431 WWL[11].n29 WWL[11].t25 260.715
R13432 WWL[11].n27 WWL[11].t23 260.715
R13433 WWL[11].n25 WWL[11].t17 260.715
R13434 WWL[11].n23 WWL[11].t26 260.715
R13435 WWL[11].n21 WWL[11].t24 260.715
R13436 WWL[11].n19 WWL[11].t12 260.715
R13437 WWL[11].n17 WWL[11].t28 260.715
R13438 WWL[11].n15 WWL[11].t15 260.715
R13439 WWL[11].n13 WWL[11].t3 260.715
R13440 WWL[11].n11 WWL[11].t29 260.715
R13441 WWL[11].n9 WWL[11].t16 260.715
R13442 WWL[11].n7 WWL[11].t5 260.715
R13443 WWL[11].n5 WWL[11].t21 260.715
R13444 WWL[11].n3 WWL[11].t11 260.715
R13445 WWL[11].n1 WWL[11].t7 260.715
R13446 WWL[11].n30 WWL[11].t27 259.254
R13447 WWL[11].n28 WWL[11].t2 259.254
R13448 WWL[11].n26 WWL[11].t13 259.254
R13449 WWL[11].n24 WWL[11].t30 259.254
R13450 WWL[11].n22 WWL[11].t20 259.254
R13451 WWL[11].n20 WWL[11].t4 259.254
R13452 WWL[11].n18 WWL[11].t18 259.254
R13453 WWL[11].n16 WWL[11].t0 259.254
R13454 WWL[11].n14 WWL[11].t22 259.254
R13455 WWL[11].n12 WWL[11].t9 259.254
R13456 WWL[11].n10 WWL[11].t31 259.254
R13457 WWL[11].n8 WWL[11].t6 259.254
R13458 WWL[11].n6 WWL[11].t8 259.254
R13459 WWL[11].n4 WWL[11].t10 259.254
R13460 WWL[11].n2 WWL[11].t1 259.254
R13461 WWL[11].n0 WWL[11].t19 259.254
R13462 WWL[11] WWL[11].n30 44.647
R13463 WWL[11].n1 WWL[11].n0 3.576
R13464 WWL[11].n3 WWL[11].n2 3.576
R13465 WWL[11].n5 WWL[11].n4 3.576
R13466 WWL[11].n7 WWL[11].n6 3.576
R13467 WWL[11].n9 WWL[11].n8 3.576
R13468 WWL[11].n11 WWL[11].n10 3.576
R13469 WWL[11].n13 WWL[11].n12 3.576
R13470 WWL[11].n15 WWL[11].n14 3.576
R13471 WWL[11].n17 WWL[11].n16 3.576
R13472 WWL[11].n19 WWL[11].n18 3.576
R13473 WWL[11].n21 WWL[11].n20 3.576
R13474 WWL[11].n23 WWL[11].n22 3.576
R13475 WWL[11].n25 WWL[11].n24 3.576
R13476 WWL[11].n27 WWL[11].n26 3.576
R13477 WWL[11].n29 WWL[11].n28 3.576
R13478 WWL[11].n2 WWL[11].n1 1.317
R13479 WWL[11].n4 WWL[11].n3 1.317
R13480 WWL[11].n6 WWL[11].n5 1.317
R13481 WWL[11].n8 WWL[11].n7 1.317
R13482 WWL[11].n10 WWL[11].n9 1.317
R13483 WWL[11].n12 WWL[11].n11 1.317
R13484 WWL[11].n14 WWL[11].n13 1.317
R13485 WWL[11].n16 WWL[11].n15 1.317
R13486 WWL[11].n18 WWL[11].n17 1.317
R13487 WWL[11].n20 WWL[11].n19 1.317
R13488 WWL[11].n22 WWL[11].n21 1.317
R13489 WWL[11].n24 WWL[11].n23 1.317
R13490 WWL[11].n26 WWL[11].n25 1.317
R13491 WWL[11].n28 WWL[11].n27 1.317
R13492 WWL[11].n30 WWL[11].n29 1.317
R13493 a_4397_975.n0 a_4397_975.t1 358.166
R13494 a_4397_975.t4 a_4397_975.t5 337.399
R13495 a_4397_975.t5 a_4397_975.t3 285.986
R13496 a_4397_975.n0 a_4397_975.t4 282.573
R13497 a_4397_975.n1 a_4397_975.t0 202.857
R13498 a_4397_975.n1 a_4397_975.n0 173.817
R13499 a_4397_975.n1 a_4397_975.t2 20.826
R13500 a_4397_975.n2 a_4397_975.n1 20.689
R13501 a_4408_n953.n25 a_4408_n953.t27 561.971
R13502 a_4408_n953.n0 a_4408_n953.t22 461.908
R13503 a_4408_n953.t8 a_4408_n953.n25 108.635
R13504 a_4408_n953.n0 a_4408_n953.t23 79.512
R13505 a_4408_n953.n24 a_4408_n953.t25 65.401
R13506 a_4408_n953.n23 a_4408_n953.t12 65.401
R13507 a_4408_n953.n22 a_4408_n953.t4 65.401
R13508 a_4408_n953.n21 a_4408_n953.t9 65.401
R13509 a_4408_n953.n20 a_4408_n953.t16 65.401
R13510 a_4408_n953.n19 a_4408_n953.t11 65.401
R13511 a_4408_n953.n18 a_4408_n953.t24 65.401
R13512 a_4408_n953.n17 a_4408_n953.t7 65.401
R13513 a_4408_n953.n16 a_4408_n953.t1 65.401
R13514 a_4408_n953.n15 a_4408_n953.t5 65.401
R13515 a_4408_n953.n14 a_4408_n953.t14 65.401
R13516 a_4408_n953.n13 a_4408_n953.t2 65.401
R13517 a_4408_n953.n12 a_4408_n953.t10 65.401
R13518 a_4408_n953.n11 a_4408_n953.t19 65.401
R13519 a_4408_n953.n10 a_4408_n953.t3 65.401
R13520 a_4408_n953.n9 a_4408_n953.t15 65.401
R13521 a_4408_n953.n8 a_4408_n953.t13 65.401
R13522 a_4408_n953.n7 a_4408_n953.t26 65.401
R13523 a_4408_n953.n6 a_4408_n953.t0 65.401
R13524 a_4408_n953.n5 a_4408_n953.t20 65.401
R13525 a_4408_n953.n4 a_4408_n953.t6 65.401
R13526 a_4408_n953.n3 a_4408_n953.t17 65.401
R13527 a_4408_n953.n2 a_4408_n953.t18 65.401
R13528 a_4408_n953.n1 a_4408_n953.t21 65.401
R13529 a_4408_n953.n1 a_4408_n953.n0 5.64
R13530 a_4408_n953.n25 a_4408_n953.n24 4.438
R13531 a_4408_n953.n23 a_4408_n953.n22 2.524
R13532 a_4408_n953.n3 a_4408_n953.n2 2.498
R13533 a_4408_n953.n17 a_4408_n953.n16 2.364
R13534 a_4408_n953.n9 a_4408_n953.n8 2.355
R13535 a_4408_n953.n2 a_4408_n953.n1 1.998
R13536 a_4408_n953.n4 a_4408_n953.n3 1.998
R13537 a_4408_n953.n5 a_4408_n953.n4 1.998
R13538 a_4408_n953.n6 a_4408_n953.n5 1.998
R13539 a_4408_n953.n7 a_4408_n953.n6 1.998
R13540 a_4408_n953.n8 a_4408_n953.n7 1.998
R13541 a_4408_n953.n10 a_4408_n953.n9 1.998
R13542 a_4408_n953.n11 a_4408_n953.n10 1.998
R13543 a_4408_n953.n12 a_4408_n953.n11 1.998
R13544 a_4408_n953.n13 a_4408_n953.n12 1.998
R13545 a_4408_n953.n14 a_4408_n953.n13 1.998
R13546 a_4408_n953.n15 a_4408_n953.n14 1.998
R13547 a_4408_n953.n16 a_4408_n953.n15 1.998
R13548 a_4408_n953.n18 a_4408_n953.n17 1.998
R13549 a_4408_n953.n19 a_4408_n953.n18 1.998
R13550 a_4408_n953.n20 a_4408_n953.n19 1.998
R13551 a_4408_n953.n21 a_4408_n953.n20 1.998
R13552 a_4408_n953.n22 a_4408_n953.n21 1.998
R13553 a_4408_n953.n24 a_4408_n953.n23 1.998
R13554 a_593_n2086.t0 a_593_n2086.t1 34.8
R13555 a_545_4887.n25 a_545_4887.t27 561.971
R13556 a_545_4887.n0 a_545_4887.t23 449.944
R13557 a_545_4887.t8 a_545_4887.n25 108.636
R13558 a_545_4887.n0 a_545_4887.t22 74.821
R13559 a_545_4887.n24 a_545_4887.t26 63.519
R13560 a_545_4887.n23 a_545_4887.t12 63.519
R13561 a_545_4887.n22 a_545_4887.t4 63.519
R13562 a_545_4887.n21 a_545_4887.t9 63.519
R13563 a_545_4887.n20 a_545_4887.t16 63.519
R13564 a_545_4887.n19 a_545_4887.t11 63.519
R13565 a_545_4887.n18 a_545_4887.t24 63.519
R13566 a_545_4887.n17 a_545_4887.t7 63.519
R13567 a_545_4887.n16 a_545_4887.t1 63.519
R13568 a_545_4887.n15 a_545_4887.t5 63.519
R13569 a_545_4887.n14 a_545_4887.t14 63.519
R13570 a_545_4887.n13 a_545_4887.t2 63.519
R13571 a_545_4887.n12 a_545_4887.t10 63.519
R13572 a_545_4887.n11 a_545_4887.t19 63.519
R13573 a_545_4887.n10 a_545_4887.t3 63.519
R13574 a_545_4887.n9 a_545_4887.t15 63.519
R13575 a_545_4887.n8 a_545_4887.t13 63.519
R13576 a_545_4887.n7 a_545_4887.t25 63.519
R13577 a_545_4887.n6 a_545_4887.t0 63.519
R13578 a_545_4887.n5 a_545_4887.t20 63.519
R13579 a_545_4887.n4 a_545_4887.t6 63.519
R13580 a_545_4887.n3 a_545_4887.t17 63.519
R13581 a_545_4887.n2 a_545_4887.t18 63.519
R13582 a_545_4887.n1 a_545_4887.t21 63.519
R13583 a_545_4887.n1 a_545_4887.n0 8.619
R13584 a_545_4887.n25 a_545_4887.n24 2.946
R13585 a_545_4887.n23 a_545_4887.n22 2.524
R13586 a_545_4887.n3 a_545_4887.n2 2.498
R13587 a_545_4887.n17 a_545_4887.n16 2.364
R13588 a_545_4887.n9 a_545_4887.n8 2.355
R13589 a_545_4887.n24 a_545_4887.n23 1.998
R13590 a_545_4887.n22 a_545_4887.n21 1.998
R13591 a_545_4887.n21 a_545_4887.n20 1.998
R13592 a_545_4887.n20 a_545_4887.n19 1.998
R13593 a_545_4887.n19 a_545_4887.n18 1.998
R13594 a_545_4887.n18 a_545_4887.n17 1.998
R13595 a_545_4887.n16 a_545_4887.n15 1.998
R13596 a_545_4887.n15 a_545_4887.n14 1.998
R13597 a_545_4887.n14 a_545_4887.n13 1.998
R13598 a_545_4887.n13 a_545_4887.n12 1.998
R13599 a_545_4887.n12 a_545_4887.n11 1.998
R13600 a_545_4887.n11 a_545_4887.n10 1.998
R13601 a_545_4887.n10 a_545_4887.n9 1.998
R13602 a_545_4887.n8 a_545_4887.n7 1.998
R13603 a_545_4887.n7 a_545_4887.n6 1.998
R13604 a_545_4887.n6 a_545_4887.n5 1.998
R13605 a_545_4887.n5 a_545_4887.n4 1.998
R13606 a_545_4887.n4 a_545_4887.n3 1.998
R13607 a_545_4887.n2 a_545_4887.n1 1.998
R13608 a_865_4445.t0 a_865_4445.t1 242.857
R13609 a_3247_3425.n0 a_3247_3425.t1 358.166
R13610 a_3247_3425.t4 a_3247_3425.t5 337.399
R13611 a_3247_3425.t5 a_3247_3425.t3 285.986
R13612 a_3247_3425.n0 a_3247_3425.t4 282.573
R13613 a_3247_3425.n1 a_3247_3425.t0 202.857
R13614 a_3247_3425.n1 a_3247_3425.n0 173.817
R13615 a_3247_3425.n1 a_3247_3425.t2 20.826
R13616 a_3247_3425.n2 a_3247_3425.n1 20.689
R13617 a_n1495_n4378.n3 a_n1495_n4378.t2 475.39
R13618 a_n1495_n4378.t5 a_n1495_n4378.t7 228.696
R13619 a_n1495_n4378.n3 a_n1495_n4378.n2 206.292
R13620 a_n1495_n4378.n2 a_n1495_n4378.t1 185.704
R13621 a_n1495_n4378.n0 a_n1495_n4378.t5 126.761
R13622 a_n1495_n4378.n1 a_n1495_n4378.t6 126.284
R13623 a_n1495_n4378.n1 a_n1495_n4378.t0 126.284
R13624 a_n1495_n4378.t3 a_n1495_n4378.n3 124.375
R13625 a_n1495_n4378.t0 a_n1495_n4378.n0 115.122
R13626 a_n1495_n4378.n0 a_n1495_n4378.t4 111.229
R13627 a_n1495_n4378.n2 a_n1495_n4378.n1 8.764
R13628 a_n1495_n5092.t0 a_n1495_n5092.t1 42.705
R13629 WWLD[7].n0 WWLD[7].t11 262.032
R13630 WWLD[7].n29 WWLD[7].t9 260.715
R13631 WWLD[7].n27 WWLD[7].t24 260.715
R13632 WWLD[7].n25 WWLD[7].t6 260.715
R13633 WWLD[7].n23 WWLD[7].t13 260.715
R13634 WWLD[7].n21 WWLD[7].t30 260.715
R13635 WWLD[7].n19 WWLD[7].t15 260.715
R13636 WWLD[7].n17 WWLD[7].t25 260.715
R13637 WWLD[7].n15 WWLD[7].t1 260.715
R13638 WWLD[7].n13 WWLD[7].t14 260.715
R13639 WWLD[7].n11 WWLD[7].t4 260.715
R13640 WWLD[7].n9 WWLD[7].t16 260.715
R13641 WWLD[7].n7 WWLD[7].t28 260.715
R13642 WWLD[7].n5 WWLD[7].t3 260.715
R13643 WWLD[7].n3 WWLD[7].t20 260.715
R13644 WWLD[7].n1 WWLD[7].t5 260.715
R13645 WWLD[7].n30 WWLD[7].t17 259.254
R13646 WWLD[7].n28 WWLD[7].t23 259.254
R13647 WWLD[7].n26 WWLD[7].t2 259.254
R13648 WWLD[7].n24 WWLD[7].t18 259.254
R13649 WWLD[7].n22 WWLD[7].t10 259.254
R13650 WWLD[7].n20 WWLD[7].t26 259.254
R13651 WWLD[7].n18 WWLD[7].t7 259.254
R13652 WWLD[7].n16 WWLD[7].t21 259.254
R13653 WWLD[7].n14 WWLD[7].t12 259.254
R13654 WWLD[7].n12 WWLD[7].t31 259.254
R13655 WWLD[7].n10 WWLD[7].t19 259.254
R13656 WWLD[7].n8 WWLD[7].t27 259.254
R13657 WWLD[7].n6 WWLD[7].t29 259.254
R13658 WWLD[7].n4 WWLD[7].t0 259.254
R13659 WWLD[7].n2 WWLD[7].t22 259.254
R13660 WWLD[7].n0 WWLD[7].t8 259.254
R13661 WWLD[7] WWLD[7].n30 44.647
R13662 WWLD[7].n1 WWLD[7].n0 3.576
R13663 WWLD[7].n3 WWLD[7].n2 3.576
R13664 WWLD[7].n5 WWLD[7].n4 3.576
R13665 WWLD[7].n7 WWLD[7].n6 3.576
R13666 WWLD[7].n9 WWLD[7].n8 3.576
R13667 WWLD[7].n11 WWLD[7].n10 3.576
R13668 WWLD[7].n13 WWLD[7].n12 3.576
R13669 WWLD[7].n15 WWLD[7].n14 3.576
R13670 WWLD[7].n17 WWLD[7].n16 3.576
R13671 WWLD[7].n19 WWLD[7].n18 3.576
R13672 WWLD[7].n21 WWLD[7].n20 3.576
R13673 WWLD[7].n23 WWLD[7].n22 3.576
R13674 WWLD[7].n25 WWLD[7].n24 3.576
R13675 WWLD[7].n27 WWLD[7].n26 3.576
R13676 WWLD[7].n29 WWLD[7].n28 3.576
R13677 WWLD[7].n2 WWLD[7].n1 1.317
R13678 WWLD[7].n4 WWLD[7].n3 1.317
R13679 WWLD[7].n6 WWLD[7].n5 1.317
R13680 WWLD[7].n8 WWLD[7].n7 1.317
R13681 WWLD[7].n10 WWLD[7].n9 1.317
R13682 WWLD[7].n12 WWLD[7].n11 1.317
R13683 WWLD[7].n14 WWLD[7].n13 1.317
R13684 WWLD[7].n16 WWLD[7].n15 1.317
R13685 WWLD[7].n18 WWLD[7].n17 1.317
R13686 WWLD[7].n20 WWLD[7].n19 1.317
R13687 WWLD[7].n22 WWLD[7].n21 1.317
R13688 WWLD[7].n24 WWLD[7].n23 1.317
R13689 WWLD[7].n26 WWLD[7].n25 1.317
R13690 WWLD[7].n28 WWLD[7].n27 1.317
R13691 WWLD[7].n30 WWLD[7].n29 1.317
R13692 a_7847_n1053.n0 a_7847_n1053.t0 358.166
R13693 a_7847_n1053.t5 a_7847_n1053.t3 337.399
R13694 a_7847_n1053.t3 a_7847_n1053.t4 285.986
R13695 a_7847_n1053.n0 a_7847_n1053.t5 282.573
R13696 a_7847_n1053.n1 a_7847_n1053.t2 202.857
R13697 a_7847_n1053.n1 a_7847_n1053.n0 173.817
R13698 a_7847_n1053.n1 a_7847_n1053.t1 20.826
R13699 a_7847_n1053.n2 a_7847_n1053.n1 20.689
R13700 a_7858_n953.n25 a_7858_n953.t27 561.971
R13701 a_7858_n953.n0 a_7858_n953.t25 461.908
R13702 a_7858_n953.t8 a_7858_n953.n25 108.635
R13703 a_7858_n953.n0 a_7858_n953.t24 79.512
R13704 a_7858_n953.n24 a_7858_n953.t14 65.401
R13705 a_7858_n953.n23 a_7858_n953.t12 65.401
R13706 a_7858_n953.n22 a_7858_n953.t4 65.401
R13707 a_7858_n953.n21 a_7858_n953.t9 65.401
R13708 a_7858_n953.n20 a_7858_n953.t17 65.401
R13709 a_7858_n953.n19 a_7858_n953.t11 65.401
R13710 a_7858_n953.n18 a_7858_n953.t23 65.401
R13711 a_7858_n953.n17 a_7858_n953.t7 65.401
R13712 a_7858_n953.n16 a_7858_n953.t1 65.401
R13713 a_7858_n953.n15 a_7858_n953.t5 65.401
R13714 a_7858_n953.n14 a_7858_n953.t15 65.401
R13715 a_7858_n953.n13 a_7858_n953.t2 65.401
R13716 a_7858_n953.n12 a_7858_n953.t10 65.401
R13717 a_7858_n953.n11 a_7858_n953.t20 65.401
R13718 a_7858_n953.n10 a_7858_n953.t3 65.401
R13719 a_7858_n953.n9 a_7858_n953.t16 65.401
R13720 a_7858_n953.n8 a_7858_n953.t13 65.401
R13721 a_7858_n953.n7 a_7858_n953.t26 65.401
R13722 a_7858_n953.n6 a_7858_n953.t0 65.401
R13723 a_7858_n953.n5 a_7858_n953.t21 65.401
R13724 a_7858_n953.n4 a_7858_n953.t6 65.401
R13725 a_7858_n953.n3 a_7858_n953.t18 65.401
R13726 a_7858_n953.n2 a_7858_n953.t19 65.401
R13727 a_7858_n953.n1 a_7858_n953.t22 65.401
R13728 a_7858_n953.n1 a_7858_n953.n0 5.64
R13729 a_7858_n953.n25 a_7858_n953.n24 4.438
R13730 a_7858_n953.n23 a_7858_n953.n22 2.524
R13731 a_7858_n953.n3 a_7858_n953.n2 2.498
R13732 a_7858_n953.n17 a_7858_n953.n16 2.364
R13733 a_7858_n953.n9 a_7858_n953.n8 2.355
R13734 a_7858_n953.n2 a_7858_n953.n1 1.998
R13735 a_7858_n953.n4 a_7858_n953.n3 1.998
R13736 a_7858_n953.n5 a_7858_n953.n4 1.998
R13737 a_7858_n953.n6 a_7858_n953.n5 1.998
R13738 a_7858_n953.n7 a_7858_n953.n6 1.998
R13739 a_7858_n953.n8 a_7858_n953.n7 1.998
R13740 a_7858_n953.n10 a_7858_n953.n9 1.998
R13741 a_7858_n953.n11 a_7858_n953.n10 1.998
R13742 a_7858_n953.n12 a_7858_n953.n11 1.998
R13743 a_7858_n953.n13 a_7858_n953.n12 1.998
R13744 a_7858_n953.n14 a_7858_n953.n13 1.998
R13745 a_7858_n953.n15 a_7858_n953.n14 1.998
R13746 a_7858_n953.n16 a_7858_n953.n15 1.998
R13747 a_7858_n953.n18 a_7858_n953.n17 1.998
R13748 a_7858_n953.n19 a_7858_n953.n18 1.998
R13749 a_7858_n953.n20 a_7858_n953.n19 1.998
R13750 a_7858_n953.n21 a_7858_n953.n20 1.998
R13751 a_7858_n953.n22 a_7858_n953.n21 1.998
R13752 a_7858_n953.n24 a_7858_n953.n23 1.998
R13753 a_7752_437.n0 a_7752_437.t1 362.857
R13754 a_7752_437.t5 a_7752_437.t4 337.399
R13755 a_7752_437.t4 a_7752_437.t3 298.839
R13756 a_7752_437.n0 a_7752_437.t5 280.405
R13757 a_7752_437.n1 a_7752_437.t2 200
R13758 a_7752_437.n1 a_7752_437.n0 172.311
R13759 a_7752_437.n2 a_7752_437.n1 24
R13760 a_7752_437.n1 a_7752_437.t0 21.212
R13761 a_7765_452.t0 a_7765_452.t1 242.857
R13762 Iref3.n0 Iref3.t5 463.921
R13763 Iref3.n14 Iref3.t4 456.275
R13764 Iref3.n13 Iref3.t13 456.275
R13765 Iref3.n12 Iref3.t6 456.275
R13766 Iref3.n11 Iref3.t12 456.275
R13767 Iref3.n10 Iref3.t11 456.275
R13768 Iref3.n9 Iref3.t15 456.275
R13769 Iref3.n8 Iref3.t2 456.275
R13770 Iref3.n7 Iref3.t9 456.275
R13771 Iref3.n6 Iref3.t1 456.275
R13772 Iref3.n5 Iref3.t8 456.275
R13773 Iref3.n4 Iref3.t0 456.275
R13774 Iref3.n3 Iref3.t7 456.275
R13775 Iref3.n2 Iref3.t10 456.275
R13776 Iref3.n1 Iref3.t3 456.275
R13777 Iref3.n0 Iref3.t14 456.275
R13778 Iref3 Iref3.n14 20.041
R13779 Iref3.n12 Iref3.n11 8.671
R13780 Iref3.n13 Iref3.n12 8.671
R13781 Iref3.n10 Iref3.n9 8.649
R13782 Iref3.n11 Iref3.n10 8.649
R13783 Iref3.n1 Iref3.n0 8.634
R13784 Iref3.n4 Iref3.n3 8.634
R13785 Iref3.n5 Iref3.n4 8.634
R13786 Iref3.n6 Iref3.n5 8.634
R13787 Iref3.n7 Iref3.n6 8.634
R13788 Iref3.n8 Iref3.n7 8.634
R13789 Iref3.n9 Iref3.n8 8.634
R13790 Iref3.n2 Iref3.n1 8.627
R13791 Iref3.n3 Iref3.n2 8.627
R13792 Iref3.n14 Iref3.n13 6.561
R13793 a_2578_n8026.t1 a_2578_n8026.t0 336.814
R13794 a_2519_n8071.t0 a_2519_n8071.t1 68.74
R13795 a_3493_n8583.n0 a_3493_n8583.t4 1465.51
R13796 a_3493_n8583.n0 a_3493_n8583.t3 712.44
R13797 a_3493_n8583.n1 a_3493_n8583.t0 375.067
R13798 a_3493_n8583.n1 a_3493_n8583.t2 272.668
R13799 a_3493_n8583.n2 a_3493_n8583.n0 143.764
R13800 a_3493_n8583.t1 a_3493_n8583.n2 78.193
R13801 a_3493_n8583.n2 a_3493_n8583.n1 4.517
R13802 a_7283_n953.n25 a_7283_n953.t27 561.971
R13803 a_7283_n953.n0 a_7283_n953.t24 461.908
R13804 a_7283_n953.t7 a_7283_n953.n25 108.635
R13805 a_7283_n953.n0 a_7283_n953.t25 79.512
R13806 a_7283_n953.n24 a_7283_n953.t13 65.401
R13807 a_7283_n953.n23 a_7283_n953.t11 65.401
R13808 a_7283_n953.n22 a_7283_n953.t3 65.401
R13809 a_7283_n953.n21 a_7283_n953.t8 65.401
R13810 a_7283_n953.n20 a_7283_n953.t19 65.401
R13811 a_7283_n953.n19 a_7283_n953.t10 65.401
R13812 a_7283_n953.n18 a_7283_n953.t23 65.401
R13813 a_7283_n953.n17 a_7283_n953.t6 65.401
R13814 a_7283_n953.n16 a_7283_n953.t1 65.401
R13815 a_7283_n953.n15 a_7283_n953.t4 65.401
R13816 a_7283_n953.n14 a_7283_n953.t14 65.401
R13817 a_7283_n953.n13 a_7283_n953.t17 65.401
R13818 a_7283_n953.n12 a_7283_n953.t9 65.401
R13819 a_7283_n953.n11 a_7283_n953.t20 65.401
R13820 a_7283_n953.n10 a_7283_n953.t2 65.401
R13821 a_7283_n953.n9 a_7283_n953.t15 65.401
R13822 a_7283_n953.n8 a_7283_n953.t12 65.401
R13823 a_7283_n953.n7 a_7283_n953.t26 65.401
R13824 a_7283_n953.n6 a_7283_n953.t0 65.401
R13825 a_7283_n953.n5 a_7283_n953.t21 65.401
R13826 a_7283_n953.n4 a_7283_n953.t5 65.401
R13827 a_7283_n953.n3 a_7283_n953.t16 65.401
R13828 a_7283_n953.n2 a_7283_n953.t18 65.401
R13829 a_7283_n953.n1 a_7283_n953.t22 65.401
R13830 a_7283_n953.n1 a_7283_n953.n0 5.64
R13831 a_7283_n953.n25 a_7283_n953.n24 4.438
R13832 a_7283_n953.n23 a_7283_n953.n22 2.524
R13833 a_7283_n953.n3 a_7283_n953.n2 2.498
R13834 a_7283_n953.n17 a_7283_n953.n16 2.364
R13835 a_7283_n953.n9 a_7283_n953.n8 2.355
R13836 a_7283_n953.n2 a_7283_n953.n1 1.998
R13837 a_7283_n953.n4 a_7283_n953.n3 1.998
R13838 a_7283_n953.n5 a_7283_n953.n4 1.998
R13839 a_7283_n953.n6 a_7283_n953.n5 1.998
R13840 a_7283_n953.n7 a_7283_n953.n6 1.998
R13841 a_7283_n953.n8 a_7283_n953.n7 1.998
R13842 a_7283_n953.n10 a_7283_n953.n9 1.998
R13843 a_7283_n953.n11 a_7283_n953.n10 1.998
R13844 a_7283_n953.n12 a_7283_n953.n11 1.998
R13845 a_7283_n953.n13 a_7283_n953.n12 1.998
R13846 a_7283_n953.n14 a_7283_n953.n13 1.998
R13847 a_7283_n953.n15 a_7283_n953.n14 1.998
R13848 a_7283_n953.n16 a_7283_n953.n15 1.998
R13849 a_7283_n953.n18 a_7283_n953.n17 1.998
R13850 a_7283_n953.n19 a_7283_n953.n18 1.998
R13851 a_7283_n953.n20 a_7283_n953.n19 1.998
R13852 a_7283_n953.n21 a_7283_n953.n20 1.998
R13853 a_7283_n953.n22 a_7283_n953.n21 1.998
R13854 a_7283_n953.n24 a_7283_n953.n23 1.998
R13855 a_7353_n2086.t0 a_7353_n2086.t1 34.8
R13856 a_2049_n4378.n3 a_2049_n4378.t2 474.093
R13857 a_2049_n4378.n3 a_2049_n4378.n2 358.637
R13858 a_2049_n4378.t5 a_2049_n4378.t7 228.696
R13859 a_2049_n4378.n2 a_2049_n4378.t1 185.704
R13860 a_2049_n4378.n0 a_2049_n4378.t5 126.761
R13861 a_2049_n4378.n1 a_2049_n4378.t6 126.284
R13862 a_2049_n4378.n1 a_2049_n4378.t0 126.284
R13863 a_2049_n4378.t0 a_2049_n4378.n0 115.122
R13864 a_2049_n4378.n0 a_2049_n4378.t4 111.229
R13865 a_2049_n4378.t3 a_2049_n4378.n3 32.938
R13866 a_2049_n4378.n2 a_2049_n4378.n1 8.764
R13867 a_4397_4445.n0 a_4397_4445.t2 358.166
R13868 a_4397_4445.t4 a_4397_4445.t5 337.399
R13869 a_4397_4445.t5 a_4397_4445.t3 285.986
R13870 a_4397_4445.n0 a_4397_4445.t4 282.573
R13871 a_4397_4445.n1 a_4397_4445.t0 202.857
R13872 a_4397_4445.n1 a_4397_4445.n0 173.817
R13873 a_4397_4445.n1 a_4397_4445.t1 20.826
R13874 a_4397_4445.n2 a_4397_4445.n1 20.689
R13875 a_4767_4445.t0 a_4767_4445.t1 242.857
R13876 a_3727_3892.n0 a_3727_3892.t2 362.857
R13877 a_3727_3892.t3 a_3727_3892.t4 337.399
R13878 a_3727_3892.t4 a_3727_3892.t5 298.839
R13879 a_3727_3892.n0 a_3727_3892.t3 280.405
R13880 a_3727_3892.n1 a_3727_3892.t0 200
R13881 a_3727_3892.n1 a_3727_3892.n0 172.311
R13882 a_3727_3892.n2 a_3727_3892.n1 24
R13883 a_3727_3892.n1 a_3727_3892.t1 21.212
R13884 a_3822_3907.n0 a_3822_3907.t2 358.166
R13885 a_3822_3907.t5 a_3822_3907.t4 337.399
R13886 a_3822_3907.t4 a_3822_3907.t3 285.986
R13887 a_3822_3907.n0 a_3822_3907.t5 282.573
R13888 a_3822_3907.n1 a_3822_3907.t0 202.857
R13889 a_3822_3907.n1 a_3822_3907.n0 173.817
R13890 a_3822_3907.n1 a_3822_3907.t1 20.826
R13891 a_3822_3907.n2 a_3822_3907.n1 20.689
R13892 a_852_437.n0 a_852_437.t1 362.857
R13893 a_852_437.t3 a_852_437.t5 337.399
R13894 a_852_437.t5 a_852_437.t4 298.839
R13895 a_852_437.n0 a_852_437.t3 280.405
R13896 a_852_437.n1 a_852_437.t2 200
R13897 a_852_437.n1 a_852_437.n0 172.311
R13898 a_852_437.n2 a_852_437.n1 24
R13899 a_852_437.n1 a_852_437.t0 21.212
R13900 a_4302_n1068.n0 a_4302_n1068.t2 362.857
R13901 a_4302_n1068.t3 a_4302_n1068.t4 337.399
R13902 a_4302_n1068.t4 a_4302_n1068.t5 298.839
R13903 a_4302_n1068.n0 a_4302_n1068.t3 280.405
R13904 a_4302_n1068.n1 a_4302_n1068.t0 200
R13905 a_4302_n1068.n1 a_4302_n1068.n0 172.311
R13906 a_4302_n1068.n2 a_4302_n1068.n1 24
R13907 a_4302_n1068.n1 a_4302_n1068.t1 21.212
R13908 a_4397_n1053.n0 a_4397_n1053.t1 358.166
R13909 a_4397_n1053.t4 a_4397_n1053.t5 337.399
R13910 a_4397_n1053.t5 a_4397_n1053.t3 285.986
R13911 a_4397_n1053.n0 a_4397_n1053.t4 282.573
R13912 a_4397_n1053.n1 a_4397_n1053.t2 202.857
R13913 a_4397_n1053.n1 a_4397_n1053.n0 173.817
R13914 a_4397_n1053.n1 a_4397_n1053.t0 20.826
R13915 a_4397_n1053.n2 a_4397_n1053.n1 20.689
R13916 a_3727_n1068.n0 a_3727_n1068.t2 362.857
R13917 a_3727_n1068.t5 a_3727_n1068.t3 337.399
R13918 a_3727_n1068.t3 a_3727_n1068.t4 298.839
R13919 a_3727_n1068.n0 a_3727_n1068.t5 280.405
R13920 a_3727_n1068.n1 a_3727_n1068.t0 200
R13921 a_3727_n1068.n1 a_3727_n1068.n0 172.311
R13922 a_3727_n1068.n2 a_3727_n1068.n1 24
R13923 a_3727_n1068.n1 a_3727_n1068.t1 21.212
R13924 a_3822_n1053.n0 a_3822_n1053.t2 358.166
R13925 a_3822_n1053.t5 a_3822_n1053.t4 337.399
R13926 a_3822_n1053.t4 a_3822_n1053.t3 285.986
R13927 a_3822_n1053.n0 a_3822_n1053.t5 282.573
R13928 a_3822_n1053.n1 a_3822_n1053.t0 202.857
R13929 a_3822_n1053.n1 a_3822_n1053.n0 173.817
R13930 a_3822_n1053.n1 a_3822_n1053.t1 20.826
R13931 a_3822_n1053.n2 a_3822_n1053.n1 20.689
R13932 a_4972_4445.n0 a_4972_4445.t0 358.166
R13933 a_4972_4445.t4 a_4972_4445.t3 337.399
R13934 a_4972_4445.t3 a_4972_4445.t5 285.986
R13935 a_4972_4445.n0 a_4972_4445.t4 282.573
R13936 a_4972_4445.n1 a_4972_4445.t1 202.857
R13937 a_4972_4445.n1 a_4972_4445.n0 173.817
R13938 a_4972_4445.n1 a_4972_4445.t2 20.826
R13939 a_4972_4445.n2 a_4972_4445.n1 20.689
R13940 a_4877_4430.n0 a_4877_4430.t2 362.857
R13941 a_4877_4430.t4 a_4877_4430.t3 337.399
R13942 a_4877_4430.t3 a_4877_4430.t5 298.839
R13943 a_4877_4430.n0 a_4877_4430.t4 280.405
R13944 a_4877_4430.n1 a_4877_4430.t0 200
R13945 a_4877_4430.n1 a_4877_4430.n0 172.311
R13946 a_4877_4430.n2 a_4877_4430.n1 24
R13947 a_4877_4430.n1 a_4877_4430.t1 21.212
R13948 a_5465_n953.t36 a_5465_n953.n46 176.385
R13949 a_5465_n953.n22 a_5465_n953.t7 67.378
R13950 a_5465_n953.n0 a_5465_n953.t5 66.92
R13951 a_5465_n953.n1 a_5465_n953.t9 66.92
R13952 a_5465_n953.n2 a_5465_n953.t12 66.92
R13953 a_5465_n953.n3 a_5465_n953.t3 66.92
R13954 a_5465_n953.n4 a_5465_n953.t1 66.92
R13955 a_5465_n953.n5 a_5465_n953.t0 66.92
R13956 a_5465_n953.n6 a_5465_n953.t42 66.92
R13957 a_5465_n953.n7 a_5465_n953.t43 66.92
R13958 a_5465_n953.n8 a_5465_n953.t25 66.92
R13959 a_5465_n953.n9 a_5465_n953.t31 66.92
R13960 a_5465_n953.n10 a_5465_n953.t19 66.92
R13961 a_5465_n953.n11 a_5465_n953.t33 66.92
R13962 a_5465_n953.n12 a_5465_n953.t29 66.92
R13963 a_5465_n953.n13 a_5465_n953.t45 66.92
R13964 a_5465_n953.n14 a_5465_n953.t48 66.92
R13965 a_5465_n953.n15 a_5465_n953.t47 66.92
R13966 a_5465_n953.n16 a_5465_n953.t18 66.92
R13967 a_5465_n953.n17 a_5465_n953.t27 66.92
R13968 a_5465_n953.n18 a_5465_n953.t22 66.92
R13969 a_5465_n953.n19 a_5465_n953.t28 66.92
R13970 a_5465_n953.n20 a_5465_n953.t4 66.92
R13971 a_5465_n953.n21 a_5465_n953.t11 66.92
R13972 a_5465_n953.n22 a_5465_n953.t16 66.92
R13973 a_5465_n953.n23 a_5465_n953.t2 65.518
R13974 a_5465_n953.n45 a_5465_n953.t13 63.519
R13975 a_5465_n953.n44 a_5465_n953.t17 63.519
R13976 a_5465_n953.n43 a_5465_n953.t8 63.519
R13977 a_5465_n953.n42 a_5465_n953.t6 63.519
R13978 a_5465_n953.n41 a_5465_n953.t37 63.519
R13979 a_5465_n953.n40 a_5465_n953.t41 63.519
R13980 a_5465_n953.n39 a_5465_n953.t21 63.519
R13981 a_5465_n953.n38 a_5465_n953.t20 63.519
R13982 a_5465_n953.n37 a_5465_n953.t23 63.519
R13983 a_5465_n953.n36 a_5465_n953.t40 63.519
R13984 a_5465_n953.n35 a_5465_n953.t32 63.519
R13985 a_5465_n953.n34 a_5465_n953.t34 63.519
R13986 a_5465_n953.n33 a_5465_n953.t38 63.519
R13987 a_5465_n953.n32 a_5465_n953.t24 63.519
R13988 a_5465_n953.n31 a_5465_n953.t44 63.519
R13989 a_5465_n953.n30 a_5465_n953.t39 63.519
R13990 a_5465_n953.n29 a_5465_n953.t35 63.519
R13991 a_5465_n953.n28 a_5465_n953.t46 63.519
R13992 a_5465_n953.n27 a_5465_n953.t30 63.519
R13993 a_5465_n953.n26 a_5465_n953.t26 63.519
R13994 a_5465_n953.n25 a_5465_n953.t10 63.519
R13995 a_5465_n953.n24 a_5465_n953.t15 63.519
R13996 a_5465_n953.n23 a_5465_n953.t14 63.519
R13997 a_5465_n953.n46 a_5465_n953.n45 18.144
R13998 a_5465_n953.n46 a_5465_n953.n0 17.125
R13999 a_5465_n953.n44 a_5465_n953.n43 2.524
R14000 a_5465_n953.n24 a_5465_n953.n23 2.498
R14001 a_5465_n953.n21 a_5465_n953.n22 2.495
R14002 a_5465_n953.n1 a_5465_n953.n2 2.459
R14003 a_5465_n953.n38 a_5465_n953.n37 2.364
R14004 a_5465_n953.n30 a_5465_n953.n29 2.355
R14005 a_5465_n953.n7 a_5465_n953.n8 2.299
R14006 a_5465_n953.n15 a_5465_n953.n16 2.29
R14007 a_5465_n953.n16 a_5465_n953.n17 2.057
R14008 a_5465_n953.n8 a_5465_n953.n9 2.057
R14009 a_5465_n953.n2 a_5465_n953.n3 2.057
R14010 a_5465_n953.n0 a_5465_n953.n1 2.057
R14011 a_5465_n953.n45 a_5465_n953.n44 1.998
R14012 a_5465_n953.n43 a_5465_n953.n42 1.998
R14013 a_5465_n953.n42 a_5465_n953.n41 1.998
R14014 a_5465_n953.n41 a_5465_n953.n40 1.998
R14015 a_5465_n953.n40 a_5465_n953.n39 1.998
R14016 a_5465_n953.n39 a_5465_n953.n38 1.998
R14017 a_5465_n953.n37 a_5465_n953.n36 1.998
R14018 a_5465_n953.n36 a_5465_n953.n35 1.998
R14019 a_5465_n953.n35 a_5465_n953.n34 1.998
R14020 a_5465_n953.n34 a_5465_n953.n33 1.998
R14021 a_5465_n953.n33 a_5465_n953.n32 1.998
R14022 a_5465_n953.n32 a_5465_n953.n31 1.998
R14023 a_5465_n953.n31 a_5465_n953.n30 1.998
R14024 a_5465_n953.n29 a_5465_n953.n28 1.998
R14025 a_5465_n953.n28 a_5465_n953.n27 1.998
R14026 a_5465_n953.n27 a_5465_n953.n26 1.998
R14027 a_5465_n953.n26 a_5465_n953.n25 1.998
R14028 a_5465_n953.n25 a_5465_n953.n24 1.998
R14029 a_5465_n953.n20 a_5465_n953.n21 1.995
R14030 a_5465_n953.n19 a_5465_n953.n20 1.995
R14031 a_5465_n953.n18 a_5465_n953.n19 1.995
R14032 a_5465_n953.n17 a_5465_n953.n18 1.995
R14033 a_5465_n953.n14 a_5465_n953.n15 1.995
R14034 a_5465_n953.n13 a_5465_n953.n14 1.995
R14035 a_5465_n953.n12 a_5465_n953.n13 1.995
R14036 a_5465_n953.n11 a_5465_n953.n12 1.995
R14037 a_5465_n953.n10 a_5465_n953.n11 1.995
R14038 a_5465_n953.n9 a_5465_n953.n10 1.995
R14039 a_5465_n953.n6 a_5465_n953.n7 1.995
R14040 a_5465_n953.n5 a_5465_n953.n6 1.995
R14041 a_5465_n953.n4 a_5465_n953.n5 1.995
R14042 a_5465_n953.n3 a_5465_n953.n4 1.995
R14043 a_5917_2180.t0 a_5917_2180.t1 242.857
R14044 a_372_693.n0 a_372_693.t1 358.166
R14045 a_372_693.t3 a_372_693.t5 337.399
R14046 a_372_693.t5 a_372_693.t4 285.986
R14047 a_372_693.n0 a_372_693.t3 282.573
R14048 a_372_693.n1 a_372_693.t0 202.857
R14049 a_372_693.n1 a_372_693.n0 173.817
R14050 a_372_693.n1 a_372_693.t2 20.826
R14051 a_372_693.n2 a_372_693.n1 20.689
R14052 a_277_678.n0 a_277_678.t1 362.857
R14053 a_277_678.t4 a_277_678.t3 337.399
R14054 a_277_678.t3 a_277_678.t5 298.839
R14055 a_277_678.n0 a_277_678.t4 280.405
R14056 a_277_678.n1 a_277_678.t2 200
R14057 a_277_678.n1 a_277_678.n0 172.311
R14058 a_277_678.n2 a_277_678.n1 24
R14059 a_277_678.n1 a_277_678.t0 21.212
R14060 a_8422_1216.n0 a_8422_1216.t2 358.166
R14061 a_8422_1216.t5 a_8422_1216.t4 337.399
R14062 a_8422_1216.t4 a_8422_1216.t3 285.986
R14063 a_8422_1216.n0 a_8422_1216.t5 282.573
R14064 a_8422_1216.n1 a_8422_1216.t1 202.857
R14065 a_8422_1216.n1 a_8422_1216.n0 173.817
R14066 a_8422_1216.n1 a_8422_1216.t0 20.826
R14067 a_8422_1216.n2 a_8422_1216.n1 20.689
R14068 a_8792_1216.t0 a_8792_1216.t1 242.857
R14069 a_6122_452.n0 a_6122_452.t1 358.166
R14070 a_6122_452.t3 a_6122_452.t5 337.399
R14071 a_6122_452.t5 a_6122_452.t4 285.986
R14072 a_6122_452.n0 a_6122_452.t3 282.573
R14073 a_6122_452.n1 a_6122_452.t0 202.857
R14074 a_6122_452.n1 a_6122_452.n0 173.817
R14075 a_6122_452.n1 a_6122_452.t2 20.826
R14076 a_6122_452.n2 a_6122_452.n1 20.689
R14077 a_6027_437.n0 a_6027_437.t1 362.857
R14078 a_6027_437.t4 a_6027_437.t3 337.399
R14079 a_6027_437.t3 a_6027_437.t5 298.839
R14080 a_6027_437.n0 a_6027_437.t4 280.405
R14081 a_6027_437.n1 a_6027_437.t2 200
R14082 a_6027_437.n1 a_6027_437.n0 172.311
R14083 a_6027_437.n2 a_6027_437.n1 24
R14084 a_6027_437.n1 a_6027_437.t0 21.212
R14085 a_7843_n2422.n3 a_7843_n2422.t2 475.39
R14086 a_7843_n2422.n3 a_7843_n2422.n2 233.133
R14087 a_7843_n2422.t5 a_7843_n2422.t7 228.696
R14088 a_7843_n2422.n2 a_7843_n2422.t1 185.704
R14089 a_7843_n2422.n0 a_7843_n2422.t5 126.761
R14090 a_7843_n2422.n1 a_7843_n2422.t6 126.284
R14091 a_7843_n2422.n1 a_7843_n2422.t0 126.284
R14092 a_7843_n2422.t3 a_7843_n2422.n3 124.375
R14093 a_7843_n2422.t0 a_7843_n2422.n0 115.122
R14094 a_7843_n2422.n0 a_7843_n2422.t4 111.229
R14095 a_7843_n2422.n2 a_7843_n2422.n1 8.764
R14096 a_11514_n5092.t0 a_11514_n5092.t1 42.705
R14097 a_9405_n7216.n0 a_9405_n7216.t4 1464.36
R14098 a_9405_n7216.n0 a_9405_n7216.t3 713.588
R14099 a_9405_n7216.n1 a_9405_n7216.t0 374.998
R14100 a_9405_n7216.n1 a_9405_n7216.t1 273.351
R14101 a_9405_n7216.n2 a_9405_n7216.n0 143.764
R14102 a_9405_n7216.t2 a_9405_n7216.n2 78.209
R14103 a_9405_n7216.n2 a_9405_n7216.n1 4.517
R14104 ADC11_OUT[2].n0 ADC11_OUT[2].t4 1354.27
R14105 ADC11_OUT[2].n0 ADC11_OUT[2].t3 821.954
R14106 ADC11_OUT[2].n3 ADC11_OUT[2].t0 339.609
R14107 ADC11_OUT[2].n2 ADC11_OUT[2].t2 266.575
R14108 ADC11_OUT[2].n1 ADC11_OUT[2].n0 149.035
R14109 ADC11_OUT[2].n1 ADC11_OUT[2].t1 46.723
R14110 ADC11_OUT[2].n3 ADC11_OUT[2].n2 44.423
R14111 ADC11_OUT[2] ADC11_OUT[2].n3 38.209
R14112 ADC11_OUT[2].n2 ADC11_OUT[2].n1 17.317
R14113 a_372_3907.n0 a_372_3907.t1 358.166
R14114 a_372_3907.t3 a_372_3907.t5 337.399
R14115 a_372_3907.t5 a_372_3907.t4 285.986
R14116 a_372_3907.n0 a_372_3907.t3 282.573
R14117 a_372_3907.n1 a_372_3907.t0 202.857
R14118 a_372_3907.n1 a_372_3907.n0 173.817
R14119 a_372_3907.n1 a_372_3907.t2 20.826
R14120 a_372_3907.n2 a_372_3907.n1 20.689
R14121 a_277_3892.n0 a_277_3892.t2 362.857
R14122 a_277_3892.t3 a_277_3892.t4 337.399
R14123 a_277_3892.t4 a_277_3892.t5 298.839
R14124 a_277_3892.n0 a_277_3892.t3 280.405
R14125 a_277_3892.n1 a_277_3892.t0 200
R14126 a_277_3892.n1 a_277_3892.n0 172.311
R14127 a_277_3892.n2 a_277_3892.n1 24
R14128 a_277_3892.n1 a_277_3892.t1 21.212
R14129 WWL[2].n0 WWL[2].t18 262.032
R14130 WWL[2].n29 WWL[2].t21 260.715
R14131 WWL[2].n27 WWL[2].t24 260.715
R14132 WWL[2].n25 WWL[2].t6 260.715
R14133 WWL[2].n23 WWL[2].t0 260.715
R14134 WWL[2].n21 WWL[2].t12 260.715
R14135 WWL[2].n19 WWL[2].t29 260.715
R14136 WWL[2].n17 WWL[2].t20 260.715
R14137 WWL[2].n15 WWL[2].t3 260.715
R14138 WWL[2].n13 WWL[2].t25 260.715
R14139 WWL[2].n11 WWL[2].t1 260.715
R14140 WWL[2].n9 WWL[2].t22 260.715
R14141 WWL[2].n7 WWL[2].t4 260.715
R14142 WWL[2].n5 WWL[2].t30 260.715
R14143 WWL[2].n3 WWL[2].t13 260.715
R14144 WWL[2].n1 WWL[2].t26 260.715
R14145 WWL[2].n30 WWL[2].t5 259.254
R14146 WWL[2].n28 WWL[2].t11 259.254
R14147 WWL[2].n26 WWL[2].t23 259.254
R14148 WWL[2].n24 WWL[2].t7 259.254
R14149 WWL[2].n22 WWL[2].t31 259.254
R14150 WWL[2].n20 WWL[2].t14 259.254
R14151 WWL[2].n18 WWL[2].t27 259.254
R14152 WWL[2].n16 WWL[2].t9 259.254
R14153 WWL[2].n14 WWL[2].t2 259.254
R14154 WWL[2].n12 WWL[2].t17 259.254
R14155 WWL[2].n10 WWL[2].t8 259.254
R14156 WWL[2].n8 WWL[2].t15 259.254
R14157 WWL[2].n6 WWL[2].t16 259.254
R14158 WWL[2].n4 WWL[2].t19 259.254
R14159 WWL[2].n2 WWL[2].t10 259.254
R14160 WWL[2].n0 WWL[2].t28 259.254
R14161 WWL[2] WWL[2].n30 44.647
R14162 WWL[2].n1 WWL[2].n0 3.576
R14163 WWL[2].n3 WWL[2].n2 3.576
R14164 WWL[2].n5 WWL[2].n4 3.576
R14165 WWL[2].n7 WWL[2].n6 3.576
R14166 WWL[2].n9 WWL[2].n8 3.576
R14167 WWL[2].n11 WWL[2].n10 3.576
R14168 WWL[2].n13 WWL[2].n12 3.576
R14169 WWL[2].n15 WWL[2].n14 3.576
R14170 WWL[2].n17 WWL[2].n16 3.576
R14171 WWL[2].n19 WWL[2].n18 3.576
R14172 WWL[2].n21 WWL[2].n20 3.576
R14173 WWL[2].n23 WWL[2].n22 3.576
R14174 WWL[2].n25 WWL[2].n24 3.576
R14175 WWL[2].n27 WWL[2].n26 3.576
R14176 WWL[2].n29 WWL[2].n28 3.576
R14177 WWL[2].n2 WWL[2].n1 1.317
R14178 WWL[2].n4 WWL[2].n3 1.317
R14179 WWL[2].n6 WWL[2].n5 1.317
R14180 WWL[2].n8 WWL[2].n7 1.317
R14181 WWL[2].n10 WWL[2].n9 1.317
R14182 WWL[2].n12 WWL[2].n11 1.317
R14183 WWL[2].n14 WWL[2].n13 1.317
R14184 WWL[2].n16 WWL[2].n15 1.317
R14185 WWL[2].n18 WWL[2].n17 1.317
R14186 WWL[2].n20 WWL[2].n19 1.317
R14187 WWL[2].n22 WWL[2].n21 1.317
R14188 WWL[2].n24 WWL[2].n23 1.317
R14189 WWL[2].n26 WWL[2].n25 1.317
R14190 WWL[2].n28 WWL[2].n27 1.317
R14191 WWL[2].n30 WWL[2].n29 1.317
R14192 a_2270_4887.n25 a_2270_4887.t27 561.971
R14193 a_2270_4887.n0 a_2270_4887.t25 449.944
R14194 a_2270_4887.t9 a_2270_4887.n25 108.636
R14195 a_2270_4887.n0 a_2270_4887.t24 74.821
R14196 a_2270_4887.n24 a_2270_4887.t15 63.519
R14197 a_2270_4887.n23 a_2270_4887.t13 63.519
R14198 a_2270_4887.n22 a_2270_4887.t4 63.519
R14199 a_2270_4887.n21 a_2270_4887.t10 63.519
R14200 a_2270_4887.n20 a_2270_4887.t18 63.519
R14201 a_2270_4887.n19 a_2270_4887.t12 63.519
R14202 a_2270_4887.n18 a_2270_4887.t26 63.519
R14203 a_2270_4887.n17 a_2270_4887.t7 63.519
R14204 a_2270_4887.n16 a_2270_4887.t3 63.519
R14205 a_2270_4887.n15 a_2270_4887.t5 63.519
R14206 a_2270_4887.n14 a_2270_4887.t16 63.519
R14207 a_2270_4887.n13 a_2270_4887.t0 63.519
R14208 a_2270_4887.n12 a_2270_4887.t11 63.519
R14209 a_2270_4887.n11 a_2270_4887.t21 63.519
R14210 a_2270_4887.n10 a_2270_4887.t8 63.519
R14211 a_2270_4887.n9 a_2270_4887.t17 63.519
R14212 a_2270_4887.n8 a_2270_4887.t14 63.519
R14213 a_2270_4887.n7 a_2270_4887.t2 63.519
R14214 a_2270_4887.n6 a_2270_4887.t1 63.519
R14215 a_2270_4887.n5 a_2270_4887.t22 63.519
R14216 a_2270_4887.n4 a_2270_4887.t6 63.519
R14217 a_2270_4887.n3 a_2270_4887.t19 63.519
R14218 a_2270_4887.n2 a_2270_4887.t20 63.519
R14219 a_2270_4887.n1 a_2270_4887.t23 63.519
R14220 a_2270_4887.n1 a_2270_4887.n0 8.619
R14221 a_2270_4887.n25 a_2270_4887.n24 2.946
R14222 a_2270_4887.n23 a_2270_4887.n22 2.524
R14223 a_2270_4887.n3 a_2270_4887.n2 2.498
R14224 a_2270_4887.n17 a_2270_4887.n16 2.364
R14225 a_2270_4887.n9 a_2270_4887.n8 2.355
R14226 a_2270_4887.n24 a_2270_4887.n23 1.998
R14227 a_2270_4887.n22 a_2270_4887.n21 1.998
R14228 a_2270_4887.n21 a_2270_4887.n20 1.998
R14229 a_2270_4887.n20 a_2270_4887.n19 1.998
R14230 a_2270_4887.n19 a_2270_4887.n18 1.998
R14231 a_2270_4887.n18 a_2270_4887.n17 1.998
R14232 a_2270_4887.n16 a_2270_4887.n15 1.998
R14233 a_2270_4887.n15 a_2270_4887.n14 1.998
R14234 a_2270_4887.n14 a_2270_4887.n13 1.998
R14235 a_2270_4887.n13 a_2270_4887.n12 1.998
R14236 a_2270_4887.n12 a_2270_4887.n11 1.998
R14237 a_2270_4887.n11 a_2270_4887.n10 1.998
R14238 a_2270_4887.n10 a_2270_4887.n9 1.998
R14239 a_2270_4887.n8 a_2270_4887.n7 1.998
R14240 a_2270_4887.n7 a_2270_4887.n6 1.998
R14241 a_2270_4887.n6 a_2270_4887.n5 1.998
R14242 a_2270_4887.n5 a_2270_4887.n4 1.998
R14243 a_2270_4887.n4 a_2270_4887.n3 1.998
R14244 a_2270_4887.n2 a_2270_4887.n1 1.998
R14245 a_2002_3169.n0 a_2002_3169.t1 362.857
R14246 a_2002_3169.t3 a_2002_3169.t5 337.399
R14247 a_2002_3169.t5 a_2002_3169.t4 298.839
R14248 a_2002_3169.n0 a_2002_3169.t3 280.405
R14249 a_2002_3169.n1 a_2002_3169.t0 200
R14250 a_2002_3169.n1 a_2002_3169.n0 172.311
R14251 a_2002_3169.n2 a_2002_3169.n1 24
R14252 a_2002_3169.n1 a_2002_3169.t2 21.212
R14253 WWL[13].n0 WWL[13].t7 262.032
R14254 WWL[13].n29 WWL[13].t19 260.715
R14255 WWL[13].n27 WWL[13].t17 260.715
R14256 WWL[13].n25 WWL[13].t11 260.715
R14257 WWL[13].n23 WWL[13].t21 260.715
R14258 WWL[13].n21 WWL[13].t18 260.715
R14259 WWL[13].n19 WWL[13].t2 260.715
R14260 WWL[13].n17 WWL[13].t22 260.715
R14261 WWL[13].n15 WWL[13].t8 260.715
R14262 WWL[13].n13 WWL[13].t27 260.715
R14263 WWL[13].n11 WWL[13].t23 260.715
R14264 WWL[13].n9 WWL[13].t9 260.715
R14265 WWL[13].n7 WWL[13].t28 260.715
R14266 WWL[13].n5 WWL[13].t16 260.715
R14267 WWL[13].n3 WWL[13].t1 260.715
R14268 WWL[13].n1 WWL[13].t29 260.715
R14269 WWL[13].n30 WWL[13].t14 259.254
R14270 WWL[13].n28 WWL[13].t6 259.254
R14271 WWL[13].n26 WWL[13].t4 259.254
R14272 WWL[13].n24 WWL[13].t25 259.254
R14273 WWL[13].n22 WWL[13].t12 259.254
R14274 WWL[13].n20 WWL[13].t30 259.254
R14275 WWL[13].n18 WWL[13].t26 259.254
R14276 WWL[13].n16 WWL[13].t15 259.254
R14277 WWL[13].n14 WWL[13].t31 259.254
R14278 WWL[13].n12 WWL[13].t20 259.254
R14279 WWL[13].n10 WWL[13].t3 259.254
R14280 WWL[13].n8 WWL[13].t0 259.254
R14281 WWL[13].n6 WWL[13].t10 259.254
R14282 WWL[13].n4 WWL[13].t5 259.254
R14283 WWL[13].n2 WWL[13].t24 259.254
R14284 WWL[13].n0 WWL[13].t13 259.254
R14285 WWL[13] WWL[13].n30 44.647
R14286 WWL[13].n1 WWL[13].n0 3.576
R14287 WWL[13].n3 WWL[13].n2 3.576
R14288 WWL[13].n5 WWL[13].n4 3.576
R14289 WWL[13].n7 WWL[13].n6 3.576
R14290 WWL[13].n9 WWL[13].n8 3.576
R14291 WWL[13].n11 WWL[13].n10 3.576
R14292 WWL[13].n13 WWL[13].n12 3.576
R14293 WWL[13].n15 WWL[13].n14 3.576
R14294 WWL[13].n17 WWL[13].n16 3.576
R14295 WWL[13].n19 WWL[13].n18 3.576
R14296 WWL[13].n21 WWL[13].n20 3.576
R14297 WWL[13].n23 WWL[13].n22 3.576
R14298 WWL[13].n25 WWL[13].n24 3.576
R14299 WWL[13].n27 WWL[13].n26 3.576
R14300 WWL[13].n29 WWL[13].n28 3.576
R14301 WWL[13].n2 WWL[13].n1 1.317
R14302 WWL[13].n4 WWL[13].n3 1.317
R14303 WWL[13].n6 WWL[13].n5 1.317
R14304 WWL[13].n8 WWL[13].n7 1.317
R14305 WWL[13].n10 WWL[13].n9 1.317
R14306 WWL[13].n12 WWL[13].n11 1.317
R14307 WWL[13].n14 WWL[13].n13 1.317
R14308 WWL[13].n16 WWL[13].n15 1.317
R14309 WWL[13].n18 WWL[13].n17 1.317
R14310 WWL[13].n20 WWL[13].n19 1.317
R14311 WWL[13].n22 WWL[13].n21 1.317
R14312 WWL[13].n24 WWL[13].n23 1.317
R14313 WWL[13].n26 WWL[13].n25 1.317
R14314 WWL[13].n28 WWL[13].n27 1.317
R14315 WWL[13].n30 WWL[13].n29 1.317
R14316 a_6697_452.n0 a_6697_452.t0 358.166
R14317 a_6697_452.t5 a_6697_452.t4 337.399
R14318 a_6697_452.t4 a_6697_452.t3 285.986
R14319 a_6697_452.n0 a_6697_452.t5 282.573
R14320 a_6697_452.n1 a_6697_452.t1 202.857
R14321 a_6697_452.n1 a_6697_452.n0 173.817
R14322 a_6697_452.n1 a_6697_452.t2 20.826
R14323 a_6697_452.n2 a_6697_452.n1 20.689
R14324 a_277_n527.n0 a_277_n527.t2 362.857
R14325 a_277_n527.t3 a_277_n527.t4 337.399
R14326 a_277_n527.t4 a_277_n527.t5 298.839
R14327 a_277_n527.n0 a_277_n527.t3 280.405
R14328 a_277_n527.n1 a_277_n527.t0 200
R14329 a_277_n527.n1 a_277_n527.n0 172.311
R14330 a_277_n527.n2 a_277_n527.n1 24
R14331 a_277_n527.n1 a_277_n527.t1 21.212
R14332 a_372_n512.n0 a_372_n512.t2 358.166
R14333 a_372_n512.t3 a_372_n512.t5 337.399
R14334 a_372_n512.t5 a_372_n512.t4 285.986
R14335 a_372_n512.n0 a_372_n512.t3 282.573
R14336 a_372_n512.n1 a_372_n512.t0 202.857
R14337 a_372_n512.n1 a_372_n512.n0 173.817
R14338 a_372_n512.n1 a_372_n512.t1 20.826
R14339 a_372_n512.n2 a_372_n512.n1 20.689
R14340 RWL[4].n0 RWL[4].t13 154.248
R14341 RWL[4].n14 RWL[4].t3 149.249
R14342 RWL[4].n13 RWL[4].t8 149.249
R14343 RWL[4].n12 RWL[4].t15 149.249
R14344 RWL[4].n11 RWL[4].t4 149.249
R14345 RWL[4].n10 RWL[4].t1 149.249
R14346 RWL[4].n9 RWL[4].t9 149.249
R14347 RWL[4].n8 RWL[4].t0 149.249
R14348 RWL[4].n7 RWL[4].t6 149.249
R14349 RWL[4].n6 RWL[4].t2 149.249
R14350 RWL[4].n5 RWL[4].t12 149.249
R14351 RWL[4].n4 RWL[4].t5 149.249
R14352 RWL[4].n3 RWL[4].t10 149.249
R14353 RWL[4].n2 RWL[4].t11 149.249
R14354 RWL[4].n1 RWL[4].t14 149.249
R14355 RWL[4].n0 RWL[4].t7 149.249
R14356 RWL[4] RWL[4].n14 42.874
R14357 RWL[4].n1 RWL[4].n0 4.999
R14358 RWL[4].n2 RWL[4].n1 4.999
R14359 RWL[4].n3 RWL[4].n2 4.999
R14360 RWL[4].n4 RWL[4].n3 4.999
R14361 RWL[4].n5 RWL[4].n4 4.999
R14362 RWL[4].n6 RWL[4].n5 4.999
R14363 RWL[4].n7 RWL[4].n6 4.999
R14364 RWL[4].n8 RWL[4].n7 4.999
R14365 RWL[4].n9 RWL[4].n8 4.999
R14366 RWL[4].n10 RWL[4].n9 4.999
R14367 RWL[4].n11 RWL[4].n10 4.999
R14368 RWL[4].n12 RWL[4].n11 4.999
R14369 RWL[4].n13 RWL[4].n12 4.999
R14370 RWL[4].n14 RWL[4].n13 4.999
R14371 a_3740_2662.t0 a_3740_2662.t1 242.857
R14372 a_8902_n1068.n0 a_8902_n1068.t1 362.857
R14373 a_8902_n1068.t4 a_8902_n1068.t5 337.399
R14374 a_8902_n1068.t5 a_8902_n1068.t3 298.839
R14375 a_8902_n1068.n0 a_8902_n1068.t4 280.405
R14376 a_8902_n1068.n1 a_8902_n1068.t2 200
R14377 a_8902_n1068.n1 a_8902_n1068.n0 172.311
R14378 a_8902_n1068.n2 a_8902_n1068.n1 24
R14379 a_8902_n1068.n1 a_8902_n1068.t0 21.212
R14380 a_3165_4148.t0 a_3165_4148.t1 242.857
R14381 a_3165_n953.t38 a_3165_n953.n46 176.385
R14382 a_3165_n953.n22 a_3165_n953.t7 67.378
R14383 a_3165_n953.n0 a_3165_n953.t12 66.92
R14384 a_3165_n953.n1 a_3165_n953.t0 66.92
R14385 a_3165_n953.n2 a_3165_n953.t4 66.92
R14386 a_3165_n953.n3 a_3165_n953.t9 66.92
R14387 a_3165_n953.n4 a_3165_n953.t21 66.92
R14388 a_3165_n953.n5 a_3165_n953.t47 66.92
R14389 a_3165_n953.n6 a_3165_n953.t42 66.92
R14390 a_3165_n953.n7 a_3165_n953.t43 66.92
R14391 a_3165_n953.n8 a_3165_n953.t24 66.92
R14392 a_3165_n953.n9 a_3165_n953.t32 66.92
R14393 a_3165_n953.n10 a_3165_n953.t17 66.92
R14394 a_3165_n953.n11 a_3165_n953.t35 66.92
R14395 a_3165_n953.n12 a_3165_n953.t30 66.92
R14396 a_3165_n953.n13 a_3165_n953.t44 66.92
R14397 a_3165_n953.n14 a_3165_n953.t46 66.92
R14398 a_3165_n953.n15 a_3165_n953.t26 66.92
R14399 a_3165_n953.n16 a_3165_n953.t16 66.92
R14400 a_3165_n953.n17 a_3165_n953.t28 66.92
R14401 a_3165_n953.n18 a_3165_n953.t20 66.92
R14402 a_3165_n953.n19 a_3165_n953.t29 66.92
R14403 a_3165_n953.n20 a_3165_n953.t3 66.92
R14404 a_3165_n953.n21 a_3165_n953.t13 66.92
R14405 a_3165_n953.n22 a_3165_n953.t15 66.92
R14406 a_3165_n953.n23 a_3165_n953.t2 65.518
R14407 a_3165_n953.n45 a_3165_n953.t8 63.519
R14408 a_3165_n953.n44 a_3165_n953.t14 63.519
R14409 a_3165_n953.n43 a_3165_n953.t6 63.519
R14410 a_3165_n953.n42 a_3165_n953.t11 63.519
R14411 a_3165_n953.n41 a_3165_n953.t34 63.519
R14412 a_3165_n953.n40 a_3165_n953.t41 63.519
R14413 a_3165_n953.n39 a_3165_n953.t19 63.519
R14414 a_3165_n953.n38 a_3165_n953.t18 63.519
R14415 a_3165_n953.n37 a_3165_n953.t22 63.519
R14416 a_3165_n953.n36 a_3165_n953.t40 63.519
R14417 a_3165_n953.n35 a_3165_n953.t33 63.519
R14418 a_3165_n953.n34 a_3165_n953.t36 63.519
R14419 a_3165_n953.n33 a_3165_n953.t25 63.519
R14420 a_3165_n953.n32 a_3165_n953.t23 63.519
R14421 a_3165_n953.n31 a_3165_n953.t48 63.519
R14422 a_3165_n953.n30 a_3165_n953.t39 63.519
R14423 a_3165_n953.n29 a_3165_n953.t37 63.519
R14424 a_3165_n953.n28 a_3165_n953.t45 63.519
R14425 a_3165_n953.n27 a_3165_n953.t31 63.519
R14426 a_3165_n953.n26 a_3165_n953.t27 63.519
R14427 a_3165_n953.n25 a_3165_n953.t5 63.519
R14428 a_3165_n953.n24 a_3165_n953.t10 63.519
R14429 a_3165_n953.n23 a_3165_n953.t1 63.519
R14430 a_3165_n953.n46 a_3165_n953.n45 18.144
R14431 a_3165_n953.n46 a_3165_n953.n0 17.125
R14432 a_3165_n953.n44 a_3165_n953.n43 2.524
R14433 a_3165_n953.n24 a_3165_n953.n23 2.498
R14434 a_3165_n953.n21 a_3165_n953.n22 2.495
R14435 a_3165_n953.n1 a_3165_n953.n2 2.459
R14436 a_3165_n953.n38 a_3165_n953.n37 2.364
R14437 a_3165_n953.n30 a_3165_n953.n29 2.355
R14438 a_3165_n953.n7 a_3165_n953.n8 2.299
R14439 a_3165_n953.n15 a_3165_n953.n16 2.29
R14440 a_3165_n953.n16 a_3165_n953.n17 2.057
R14441 a_3165_n953.n8 a_3165_n953.n9 2.057
R14442 a_3165_n953.n2 a_3165_n953.n3 2.057
R14443 a_3165_n953.n0 a_3165_n953.n1 2.057
R14444 a_3165_n953.n45 a_3165_n953.n44 1.998
R14445 a_3165_n953.n43 a_3165_n953.n42 1.998
R14446 a_3165_n953.n42 a_3165_n953.n41 1.998
R14447 a_3165_n953.n41 a_3165_n953.n40 1.998
R14448 a_3165_n953.n40 a_3165_n953.n39 1.998
R14449 a_3165_n953.n39 a_3165_n953.n38 1.998
R14450 a_3165_n953.n37 a_3165_n953.n36 1.998
R14451 a_3165_n953.n36 a_3165_n953.n35 1.998
R14452 a_3165_n953.n35 a_3165_n953.n34 1.998
R14453 a_3165_n953.n34 a_3165_n953.n33 1.998
R14454 a_3165_n953.n33 a_3165_n953.n32 1.998
R14455 a_3165_n953.n32 a_3165_n953.n31 1.998
R14456 a_3165_n953.n31 a_3165_n953.n30 1.998
R14457 a_3165_n953.n29 a_3165_n953.n28 1.998
R14458 a_3165_n953.n28 a_3165_n953.n27 1.998
R14459 a_3165_n953.n27 a_3165_n953.n26 1.998
R14460 a_3165_n953.n26 a_3165_n953.n25 1.998
R14461 a_3165_n953.n25 a_3165_n953.n24 1.998
R14462 a_3165_n953.n20 a_3165_n953.n21 1.995
R14463 a_3165_n953.n19 a_3165_n953.n20 1.995
R14464 a_3165_n953.n18 a_3165_n953.n19 1.995
R14465 a_3165_n953.n17 a_3165_n953.n18 1.995
R14466 a_3165_n953.n14 a_3165_n953.n15 1.995
R14467 a_3165_n953.n13 a_3165_n953.n14 1.995
R14468 a_3165_n953.n12 a_3165_n953.n13 1.995
R14469 a_3165_n953.n11 a_3165_n953.n12 1.995
R14470 a_3165_n953.n10 a_3165_n953.n11 1.995
R14471 a_3165_n953.n9 a_3165_n953.n10 1.995
R14472 a_3165_n953.n6 a_3165_n953.n7 1.995
R14473 a_3165_n953.n5 a_3165_n953.n6 1.995
R14474 a_3165_n953.n4 a_3165_n953.n5 1.995
R14475 a_3165_n953.n3 a_3165_n953.n4 1.995
R14476 a_6027_4133.n0 a_6027_4133.t2 362.857
R14477 a_6027_4133.t5 a_6027_4133.t3 337.399
R14478 a_6027_4133.t3 a_6027_4133.t4 298.839
R14479 a_6027_4133.n0 a_6027_4133.t5 280.405
R14480 a_6027_4133.n1 a_6027_4133.t0 200
R14481 a_6027_4133.n1 a_6027_4133.n0 172.311
R14482 a_6027_4133.n2 a_6027_4133.n1 24
R14483 a_6027_4133.n1 a_6027_4133.t1 21.212
R14484 a_6122_4148.n0 a_6122_4148.t1 358.166
R14485 a_6122_4148.t4 a_6122_4148.t3 337.399
R14486 a_6122_4148.t3 a_6122_4148.t5 285.986
R14487 a_6122_4148.n0 a_6122_4148.t4 282.573
R14488 a_6122_4148.n1 a_6122_4148.t2 202.857
R14489 a_6122_4148.n1 a_6122_4148.n0 173.817
R14490 a_6122_4148.n1 a_6122_4148.t0 20.826
R14491 a_6122_4148.n2 a_6122_4148.n1 20.689
R14492 a_6040_3184.t0 a_6040_3184.t1 242.857
R14493 a_7177_2165.n0 a_7177_2165.t1 362.857
R14494 a_7177_2165.t5 a_7177_2165.t3 337.399
R14495 a_7177_2165.t3 a_7177_2165.t4 298.839
R14496 a_7177_2165.n0 a_7177_2165.t5 280.405
R14497 a_7177_2165.n1 a_7177_2165.t0 200
R14498 a_7177_2165.n1 a_7177_2165.n0 172.311
R14499 a_7177_2165.n2 a_7177_2165.n1 24
R14500 a_7177_2165.n1 a_7177_2165.t2 21.212
R14501 a_7272_2180.n0 a_7272_2180.t1 358.166
R14502 a_7272_2180.t3 a_7272_2180.t5 337.399
R14503 a_7272_2180.t5 a_7272_2180.t4 285.986
R14504 a_7272_2180.n0 a_7272_2180.t3 282.573
R14505 a_7272_2180.n1 a_7272_2180.t2 202.857
R14506 a_7272_2180.n1 a_7272_2180.n0 173.817
R14507 a_7272_2180.n1 a_7272_2180.t0 20.826
R14508 a_7272_2180.n2 a_7272_2180.n1 20.689
R14509 a_2002_1683.n0 a_2002_1683.t1 362.857
R14510 a_2002_1683.t3 a_2002_1683.t5 337.399
R14511 a_2002_1683.t5 a_2002_1683.t4 298.839
R14512 a_2002_1683.n0 a_2002_1683.t3 280.405
R14513 a_2002_1683.n1 a_2002_1683.t0 200
R14514 a_2002_1683.n1 a_2002_1683.n0 172.311
R14515 a_2002_1683.n2 a_2002_1683.n1 24
R14516 a_2002_1683.n1 a_2002_1683.t2 21.212
R14517 a_2097_1698.n0 a_2097_1698.t1 358.166
R14518 a_2097_1698.t5 a_2097_1698.t3 337.399
R14519 a_2097_1698.t3 a_2097_1698.t4 285.986
R14520 a_2097_1698.n0 a_2097_1698.t5 282.573
R14521 a_2097_1698.n1 a_2097_1698.t2 202.857
R14522 a_2097_1698.n1 a_2097_1698.n0 173.817
R14523 a_2097_1698.n1 a_2097_1698.t0 20.826
R14524 a_2097_1698.n2 a_2097_1698.n1 20.689
R14525 a_1892_n512.t0 a_1892_n512.t1 242.857
R14526 a_8997_n30.n0 a_8997_n30.t2 358.166
R14527 a_8997_n30.t4 a_8997_n30.t3 337.399
R14528 a_8997_n30.t3 a_8997_n30.t5 285.986
R14529 a_8997_n30.n0 a_8997_n30.t4 282.573
R14530 a_8997_n30.n1 a_8997_n30.t0 202.857
R14531 a_8997_n30.n1 a_8997_n30.n0 173.817
R14532 a_8997_n30.n1 a_8997_n30.t1 20.826
R14533 a_8997_n30.n2 a_8997_n30.n1 20.689
R14534 a_8902_n45.n0 a_8902_n45.t1 362.857
R14535 a_8902_n45.t5 a_8902_n45.t4 337.399
R14536 a_8902_n45.t4 a_8902_n45.t3 298.839
R14537 a_8902_n45.n0 a_8902_n45.t5 280.405
R14538 a_8902_n45.n1 a_8902_n45.t2 200
R14539 a_8902_n45.n1 a_8902_n45.n0 172.311
R14540 a_8902_n45.n2 a_8902_n45.n1 24
R14541 a_8902_n45.n1 a_8902_n45.t0 21.212
R14542 a_7272_3907.n0 a_7272_3907.t1 358.166
R14543 a_7272_3907.t3 a_7272_3907.t5 337.399
R14544 a_7272_3907.t5 a_7272_3907.t4 285.986
R14545 a_7272_3907.n0 a_7272_3907.t3 282.573
R14546 a_7272_3907.n1 a_7272_3907.t0 202.857
R14547 a_7272_3907.n1 a_7272_3907.n0 173.817
R14548 a_7272_3907.n1 a_7272_3907.t2 20.826
R14549 a_7272_3907.n2 a_7272_3907.n1 20.689
R14550 a_7847_1457.n0 a_7847_1457.t0 358.166
R14551 a_7847_1457.t5 a_7847_1457.t3 337.399
R14552 a_7847_1457.t3 a_7847_1457.t4 285.986
R14553 a_7847_1457.n0 a_7847_1457.t5 282.573
R14554 a_7847_1457.n1 a_7847_1457.t1 202.857
R14555 a_7847_1457.n1 a_7847_1457.n0 173.817
R14556 a_7847_1457.n1 a_7847_1457.t2 20.826
R14557 a_7847_1457.n2 a_7847_1457.n1 20.689
R14558 a_13637_n6503.n0 a_13637_n6503.t1 65.064
R14559 a_13637_n6503.t0 a_13637_n6503.n0 42.011
R14560 a_13637_n6503.n0 a_13637_n6503.t2 2.113
R14561 RWLB[5].n0 RWLB[5].t14 154.228
R14562 RWLB[5].n14 RWLB[5].t15 149.249
R14563 RWLB[5].n13 RWLB[5].t1 149.249
R14564 RWLB[5].n12 RWLB[5].t12 149.249
R14565 RWLB[5].n11 RWLB[5].t6 149.249
R14566 RWLB[5].n10 RWLB[5].t0 149.249
R14567 RWLB[5].n9 RWLB[5].t3 149.249
R14568 RWLB[5].n8 RWLB[5].t4 149.249
R14569 RWLB[5].n7 RWLB[5].t9 149.249
R14570 RWLB[5].n6 RWLB[5].t2 149.249
R14571 RWLB[5].n5 RWLB[5].t7 149.249
R14572 RWLB[5].n4 RWLB[5].t8 149.249
R14573 RWLB[5].n3 RWLB[5].t13 149.249
R14574 RWLB[5].n2 RWLB[5].t5 149.249
R14575 RWLB[5].n1 RWLB[5].t11 149.249
R14576 RWLB[5].n0 RWLB[5].t10 149.249
R14577 RWLB[5] RWLB[5].n14 47.816
R14578 RWLB[5].n1 RWLB[5].n0 4.979
R14579 RWLB[5].n2 RWLB[5].n1 4.979
R14580 RWLB[5].n3 RWLB[5].n2 4.979
R14581 RWLB[5].n4 RWLB[5].n3 4.979
R14582 RWLB[5].n5 RWLB[5].n4 4.979
R14583 RWLB[5].n6 RWLB[5].n5 4.979
R14584 RWLB[5].n7 RWLB[5].n6 4.979
R14585 RWLB[5].n8 RWLB[5].n7 4.979
R14586 RWLB[5].n9 RWLB[5].n8 4.979
R14587 RWLB[5].n10 RWLB[5].n9 4.979
R14588 RWLB[5].n11 RWLB[5].n10 4.979
R14589 RWLB[5].n12 RWLB[5].n11 4.979
R14590 RWLB[5].n13 RWLB[5].n12 4.979
R14591 RWLB[5].n14 RWLB[5].n13 4.979
R14592 a_3042_2421.t0 a_3042_2421.t1 242.857
R14593 a_6027_960.n0 a_6027_960.t1 362.857
R14594 a_6027_960.t3 a_6027_960.t5 337.399
R14595 a_6027_960.t5 a_6027_960.t4 298.839
R14596 a_6027_960.n0 a_6027_960.t3 280.405
R14597 a_6027_960.n1 a_6027_960.t0 200
R14598 a_6027_960.n1 a_6027_960.n0 172.311
R14599 a_6027_960.n2 a_6027_960.n1 24
R14600 a_6027_960.n1 a_6027_960.t2 21.212
R14601 a_6122_975.n0 a_6122_975.t2 358.166
R14602 a_6122_975.t3 a_6122_975.t5 337.399
R14603 a_6122_975.t5 a_6122_975.t4 285.986
R14604 a_6122_975.n0 a_6122_975.t3 282.573
R14605 a_6122_975.n1 a_6122_975.t0 202.857
R14606 a_6122_975.n1 a_6122_975.n0 173.817
R14607 a_6122_975.n1 a_6122_975.t1 20.826
R14608 a_6122_975.n2 a_6122_975.n1 20.689
R14609 a_1120_4887.n25 a_1120_4887.t27 561.971
R14610 a_1120_4887.n0 a_1120_4887.t26 449.944
R14611 a_1120_4887.t8 a_1120_4887.n25 108.636
R14612 a_1120_4887.n0 a_1120_4887.t25 74.821
R14613 a_1120_4887.n24 a_1120_4887.t15 63.519
R14614 a_1120_4887.n23 a_1120_4887.t13 63.519
R14615 a_1120_4887.n22 a_1120_4887.t4 63.519
R14616 a_1120_4887.n21 a_1120_4887.t9 63.519
R14617 a_1120_4887.n20 a_1120_4887.t18 63.519
R14618 a_1120_4887.n19 a_1120_4887.t11 63.519
R14619 a_1120_4887.n18 a_1120_4887.t12 63.519
R14620 a_1120_4887.n17 a_1120_4887.t7 63.519
R14621 a_1120_4887.n16 a_1120_4887.t2 63.519
R14622 a_1120_4887.n15 a_1120_4887.t5 63.519
R14623 a_1120_4887.n14 a_1120_4887.t16 63.519
R14624 a_1120_4887.n13 a_1120_4887.t19 63.519
R14625 a_1120_4887.n12 a_1120_4887.t10 63.519
R14626 a_1120_4887.n11 a_1120_4887.t22 63.519
R14627 a_1120_4887.n10 a_1120_4887.t3 63.519
R14628 a_1120_4887.n9 a_1120_4887.t17 63.519
R14629 a_1120_4887.n8 a_1120_4887.t14 63.519
R14630 a_1120_4887.n7 a_1120_4887.t1 63.519
R14631 a_1120_4887.n6 a_1120_4887.t0 63.519
R14632 a_1120_4887.n5 a_1120_4887.t23 63.519
R14633 a_1120_4887.n4 a_1120_4887.t6 63.519
R14634 a_1120_4887.n3 a_1120_4887.t20 63.519
R14635 a_1120_4887.n2 a_1120_4887.t21 63.519
R14636 a_1120_4887.n1 a_1120_4887.t24 63.519
R14637 a_1120_4887.n1 a_1120_4887.n0 8.619
R14638 a_1120_4887.n25 a_1120_4887.n24 2.946
R14639 a_1120_4887.n23 a_1120_4887.n22 2.524
R14640 a_1120_4887.n3 a_1120_4887.n2 2.498
R14641 a_1120_4887.n17 a_1120_4887.n16 2.364
R14642 a_1120_4887.n9 a_1120_4887.n8 2.355
R14643 a_1120_4887.n24 a_1120_4887.n23 1.998
R14644 a_1120_4887.n22 a_1120_4887.n21 1.998
R14645 a_1120_4887.n21 a_1120_4887.n20 1.998
R14646 a_1120_4887.n20 a_1120_4887.n19 1.998
R14647 a_1120_4887.n19 a_1120_4887.n18 1.998
R14648 a_1120_4887.n18 a_1120_4887.n17 1.998
R14649 a_1120_4887.n16 a_1120_4887.n15 1.998
R14650 a_1120_4887.n15 a_1120_4887.n14 1.998
R14651 a_1120_4887.n14 a_1120_4887.n13 1.998
R14652 a_1120_4887.n13 a_1120_4887.n12 1.998
R14653 a_1120_4887.n12 a_1120_4887.n11 1.998
R14654 a_1120_4887.n11 a_1120_4887.n10 1.998
R14655 a_1120_4887.n10 a_1120_4887.n9 1.998
R14656 a_1120_4887.n8 a_1120_4887.n7 1.998
R14657 a_1120_4887.n7 a_1120_4887.n6 1.998
R14658 a_1120_4887.n6 a_1120_4887.n5 1.998
R14659 a_1120_4887.n5 a_1120_4887.n4 1.998
R14660 a_1120_4887.n4 a_1120_4887.n3 1.998
R14661 a_1120_4887.n2 a_1120_4887.n1 1.998
R14662 a_852_678.n0 a_852_678.t2 362.857
R14663 a_852_678.t4 a_852_678.t3 337.399
R14664 a_852_678.t3 a_852_678.t5 298.839
R14665 a_852_678.n0 a_852_678.t4 280.405
R14666 a_852_678.n1 a_852_678.t0 200
R14667 a_852_678.n1 a_852_678.n0 172.311
R14668 a_852_678.n2 a_852_678.n1 24
R14669 a_852_678.n1 a_852_678.t1 21.212
R14670 RWL[12].n0 RWL[12].t10 154.248
R14671 RWL[12].n14 RWL[12].t7 149.249
R14672 RWL[12].n13 RWL[12].t4 149.249
R14673 RWL[12].n12 RWL[12].t2 149.249
R14674 RWL[12].n11 RWL[12].t12 149.249
R14675 RWL[12].n10 RWL[12].t6 149.249
R14676 RWL[12].n9 RWL[12].t14 149.249
R14677 RWL[12].n8 RWL[12].t13 149.249
R14678 RWL[12].n7 RWL[12].t8 149.249
R14679 RWL[12].n6 RWL[12].t15 149.249
R14680 RWL[12].n5 RWL[12].t9 149.249
R14681 RWL[12].n4 RWL[12].t1 149.249
R14682 RWL[12].n3 RWL[12].t0 149.249
R14683 RWL[12].n2 RWL[12].t5 149.249
R14684 RWL[12].n1 RWL[12].t3 149.249
R14685 RWL[12].n0 RWL[12].t11 149.249
R14686 RWL[12] RWL[12].n14 42.874
R14687 RWL[12].n1 RWL[12].n0 4.999
R14688 RWL[12].n2 RWL[12].n1 4.999
R14689 RWL[12].n3 RWL[12].n2 4.999
R14690 RWL[12].n4 RWL[12].n3 4.999
R14691 RWL[12].n5 RWL[12].n4 4.999
R14692 RWL[12].n6 RWL[12].n5 4.999
R14693 RWL[12].n7 RWL[12].n6 4.999
R14694 RWL[12].n8 RWL[12].n7 4.999
R14695 RWL[12].n9 RWL[12].n8 4.999
R14696 RWL[12].n10 RWL[12].n9 4.999
R14697 RWL[12].n11 RWL[12].n10 4.999
R14698 RWL[12].n12 RWL[12].n11 4.999
R14699 RWL[12].n13 RWL[12].n12 4.999
R14700 RWL[12].n14 RWL[12].n13 4.999
R14701 a_6615_693.t0 a_6615_693.t1 242.857
R14702 a_6615_n953.t42 a_6615_n953.n46 176.385
R14703 a_6615_n953.n22 a_6615_n953.t2 67.378
R14704 a_6615_n953.n0 a_6615_n953.t7 66.92
R14705 a_6615_n953.n1 a_6615_n953.t10 66.92
R14706 a_6615_n953.n2 a_6615_n953.t8 66.92
R14707 a_6615_n953.n3 a_6615_n953.t3 66.92
R14708 a_6615_n953.n4 a_6615_n953.t23 66.92
R14709 a_6615_n953.n5 a_6615_n953.t48 66.92
R14710 a_6615_n953.n6 a_6615_n953.t44 66.92
R14711 a_6615_n953.n7 a_6615_n953.t31 66.92
R14712 a_6615_n953.n8 a_6615_n953.t26 66.92
R14713 a_6615_n953.n9 a_6615_n953.t35 66.92
R14714 a_6615_n953.n10 a_6615_n953.t18 66.92
R14715 a_6615_n953.n11 a_6615_n953.t37 66.92
R14716 a_6615_n953.n12 a_6615_n953.t32 66.92
R14717 a_6615_n953.n13 a_6615_n953.t45 66.92
R14718 a_6615_n953.n14 a_6615_n953.t47 66.92
R14719 a_6615_n953.n15 a_6615_n953.t27 66.92
R14720 a_6615_n953.n16 a_6615_n953.t17 66.92
R14721 a_6615_n953.n17 a_6615_n953.t28 66.92
R14722 a_6615_n953.n18 a_6615_n953.t21 66.92
R14723 a_6615_n953.n19 a_6615_n953.t29 66.92
R14724 a_6615_n953.n20 a_6615_n953.t4 66.92
R14725 a_6615_n953.n21 a_6615_n953.t16 66.92
R14726 a_6615_n953.n22 a_6615_n953.t5 66.92
R14727 a_6615_n953.n23 a_6615_n953.t9 65.518
R14728 a_6615_n953.n45 a_6615_n953.t13 63.519
R14729 a_6615_n953.n44 a_6615_n953.t14 63.519
R14730 a_6615_n953.n43 a_6615_n953.t12 63.519
R14731 a_6615_n953.n42 a_6615_n953.t11 63.519
R14732 a_6615_n953.n41 a_6615_n953.t39 63.519
R14733 a_6615_n953.n40 a_6615_n953.t43 63.519
R14734 a_6615_n953.n39 a_6615_n953.t20 63.519
R14735 a_6615_n953.n38 a_6615_n953.t19 63.519
R14736 a_6615_n953.n37 a_6615_n953.t24 63.519
R14737 a_6615_n953.n36 a_6615_n953.t41 63.519
R14738 a_6615_n953.n35 a_6615_n953.t36 63.519
R14739 a_6615_n953.n34 a_6615_n953.t34 63.519
R14740 a_6615_n953.n33 a_6615_n953.t0 63.519
R14741 a_6615_n953.n32 a_6615_n953.t25 63.519
R14742 a_6615_n953.n31 a_6615_n953.t22 63.519
R14743 a_6615_n953.n30 a_6615_n953.t40 63.519
R14744 a_6615_n953.n29 a_6615_n953.t38 63.519
R14745 a_6615_n953.n28 a_6615_n953.t46 63.519
R14746 a_6615_n953.n27 a_6615_n953.t33 63.519
R14747 a_6615_n953.n26 a_6615_n953.t30 63.519
R14748 a_6615_n953.n25 a_6615_n953.t6 63.519
R14749 a_6615_n953.n24 a_6615_n953.t15 63.519
R14750 a_6615_n953.n23 a_6615_n953.t1 63.519
R14751 a_6615_n953.n46 a_6615_n953.n45 18.144
R14752 a_6615_n953.n46 a_6615_n953.n0 17.125
R14753 a_6615_n953.n44 a_6615_n953.n43 2.524
R14754 a_6615_n953.n24 a_6615_n953.n23 2.498
R14755 a_6615_n953.n21 a_6615_n953.n22 2.495
R14756 a_6615_n953.n1 a_6615_n953.n2 2.459
R14757 a_6615_n953.n38 a_6615_n953.n37 2.364
R14758 a_6615_n953.n30 a_6615_n953.n29 2.355
R14759 a_6615_n953.n7 a_6615_n953.n8 2.299
R14760 a_6615_n953.n15 a_6615_n953.n16 2.29
R14761 a_6615_n953.n16 a_6615_n953.n17 2.057
R14762 a_6615_n953.n8 a_6615_n953.n9 2.057
R14763 a_6615_n953.n2 a_6615_n953.n3 2.057
R14764 a_6615_n953.n0 a_6615_n953.n1 2.057
R14765 a_6615_n953.n45 a_6615_n953.n44 1.998
R14766 a_6615_n953.n43 a_6615_n953.n42 1.998
R14767 a_6615_n953.n42 a_6615_n953.n41 1.998
R14768 a_6615_n953.n41 a_6615_n953.n40 1.998
R14769 a_6615_n953.n40 a_6615_n953.n39 1.998
R14770 a_6615_n953.n39 a_6615_n953.n38 1.998
R14771 a_6615_n953.n37 a_6615_n953.n36 1.998
R14772 a_6615_n953.n36 a_6615_n953.n35 1.998
R14773 a_6615_n953.n35 a_6615_n953.n34 1.998
R14774 a_6615_n953.n34 a_6615_n953.n33 1.998
R14775 a_6615_n953.n33 a_6615_n953.n32 1.998
R14776 a_6615_n953.n32 a_6615_n953.n31 1.998
R14777 a_6615_n953.n31 a_6615_n953.n30 1.998
R14778 a_6615_n953.n29 a_6615_n953.n28 1.998
R14779 a_6615_n953.n28 a_6615_n953.n27 1.998
R14780 a_6615_n953.n27 a_6615_n953.n26 1.998
R14781 a_6615_n953.n26 a_6615_n953.n25 1.998
R14782 a_6615_n953.n25 a_6615_n953.n24 1.998
R14783 a_6615_n953.n20 a_6615_n953.n21 1.995
R14784 a_6615_n953.n19 a_6615_n953.n20 1.995
R14785 a_6615_n953.n18 a_6615_n953.n19 1.995
R14786 a_6615_n953.n17 a_6615_n953.n18 1.995
R14787 a_6615_n953.n14 a_6615_n953.n15 1.995
R14788 a_6615_n953.n13 a_6615_n953.n14 1.995
R14789 a_6615_n953.n12 a_6615_n953.n13 1.995
R14790 a_6615_n953.n11 a_6615_n953.n12 1.995
R14791 a_6615_n953.n10 a_6615_n953.n11 1.995
R14792 a_6615_n953.n9 a_6615_n953.n10 1.995
R14793 a_6615_n953.n6 a_6615_n953.n7 1.995
R14794 a_6615_n953.n5 a_6615_n953.n6 1.995
R14795 a_6615_n953.n4 a_6615_n953.n5 1.995
R14796 a_6615_n953.n3 a_6615_n953.n4 1.995
R14797 a_6697_n512.n0 a_6697_n512.t1 358.166
R14798 a_6697_n512.t3 a_6697_n512.t4 337.399
R14799 a_6697_n512.t4 a_6697_n512.t5 285.986
R14800 a_6697_n512.n0 a_6697_n512.t3 282.573
R14801 a_6697_n512.n1 a_6697_n512.t0 202.857
R14802 a_6697_n512.n1 a_6697_n512.n0 173.817
R14803 a_6697_n512.n1 a_6697_n512.t2 20.826
R14804 a_6697_n512.n2 a_6697_n512.n1 20.689
R14805 a_6602_n527.n0 a_6602_n527.t2 362.857
R14806 a_6602_n527.t3 a_6602_n527.t5 337.399
R14807 a_6602_n527.t5 a_6602_n527.t4 298.839
R14808 a_6602_n527.n0 a_6602_n527.t3 280.405
R14809 a_6602_n527.n1 a_6602_n527.t0 200
R14810 a_6602_n527.n1 a_6602_n527.n0 172.311
R14811 a_6602_n527.n2 a_6602_n527.n1 24
R14812 a_6602_n527.n1 a_6602_n527.t1 21.212
R14813 a_2097_3184.n0 a_2097_3184.t2 358.166
R14814 a_2097_3184.t4 a_2097_3184.t5 337.399
R14815 a_2097_3184.t5 a_2097_3184.t3 285.986
R14816 a_2097_3184.n0 a_2097_3184.t4 282.573
R14817 a_2097_3184.n1 a_2097_3184.t0 202.857
R14818 a_2097_3184.n1 a_2097_3184.n0 173.817
R14819 a_2097_3184.n1 a_2097_3184.t1 20.826
R14820 a_2097_3184.n2 a_2097_3184.n1 20.689
R14821 a_2467_3184.t0 a_2467_3184.t1 242.857
R14822 a_3042_n271.t0 a_3042_n271.t1 242.857
R14823 a_3227_n2234.n2 a_3227_n2234.t0 282.97
R14824 a_3227_n2234.n1 a_3227_n2234.t2 240.683
R14825 a_3227_n2234.n0 a_3227_n2234.t3 209.208
R14826 a_3227_n2234.n0 a_3227_n2234.t4 194.167
R14827 a_3227_n2234.t1 a_3227_n2234.n2 183.404
R14828 a_3227_n2234.n1 a_3227_n2234.n0 14.805
R14829 a_3227_n2234.n2 a_3227_n2234.n1 6.415
R14830 a_3468_n2086.t0 a_3468_n2086.t1 34.8
R14831 a_5547_693.n0 a_5547_693.t1 358.166
R14832 a_5547_693.t4 a_5547_693.t3 337.399
R14833 a_5547_693.t3 a_5547_693.t5 285.986
R14834 a_5547_693.n0 a_5547_693.t4 282.573
R14835 a_5547_693.n1 a_5547_693.t0 202.857
R14836 a_5547_693.n1 a_5547_693.n0 173.817
R14837 a_5547_693.n1 a_5547_693.t2 20.826
R14838 a_5547_693.n2 a_5547_693.n1 20.689
R14839 a_5452_678.n0 a_5452_678.t1 362.857
R14840 a_5452_678.t4 a_5452_678.t3 337.399
R14841 a_5452_678.t3 a_5452_678.t5 298.839
R14842 a_5452_678.n0 a_5452_678.t4 280.405
R14843 a_5452_678.n1 a_5452_678.t2 200
R14844 a_5452_678.n1 a_5452_678.n0 172.311
R14845 a_5452_678.n2 a_5452_678.n1 24
R14846 a_5452_678.n1 a_5452_678.t0 21.212
R14847 WWLD[0].n0 WWLD[0].t0 262.032
R14848 WWLD[0].n29 WWLD[0].t3 260.715
R14849 WWLD[0].n27 WWLD[0].t6 260.715
R14850 WWLD[0].n25 WWLD[0].t20 260.715
R14851 WWLD[0].n23 WWLD[0].t14 260.715
R14852 WWLD[0].n21 WWLD[0].t26 260.715
R14853 WWLD[0].n19 WWLD[0].t11 260.715
R14854 WWLD[0].n17 WWLD[0].t2 260.715
R14855 WWLD[0].n15 WWLD[0].t17 260.715
R14856 WWLD[0].n13 WWLD[0].t7 260.715
R14857 WWLD[0].n11 WWLD[0].t15 260.715
R14858 WWLD[0].n9 WWLD[0].t4 260.715
R14859 WWLD[0].n7 WWLD[0].t18 260.715
R14860 WWLD[0].n5 WWLD[0].t12 260.715
R14861 WWLD[0].n3 WWLD[0].t27 260.715
R14862 WWLD[0].n1 WWLD[0].t8 260.715
R14863 WWLD[0].n30 WWLD[0].t19 259.254
R14864 WWLD[0].n28 WWLD[0].t25 259.254
R14865 WWLD[0].n26 WWLD[0].t5 259.254
R14866 WWLD[0].n24 WWLD[0].t21 259.254
R14867 WWLD[0].n22 WWLD[0].t13 259.254
R14868 WWLD[0].n20 WWLD[0].t28 259.254
R14869 WWLD[0].n18 WWLD[0].t9 259.254
R14870 WWLD[0].n16 WWLD[0].t23 259.254
R14871 WWLD[0].n14 WWLD[0].t16 259.254
R14872 WWLD[0].n12 WWLD[0].t31 259.254
R14873 WWLD[0].n10 WWLD[0].t22 259.254
R14874 WWLD[0].n8 WWLD[0].t29 259.254
R14875 WWLD[0].n6 WWLD[0].t30 259.254
R14876 WWLD[0].n4 WWLD[0].t1 259.254
R14877 WWLD[0].n2 WWLD[0].t24 259.254
R14878 WWLD[0].n0 WWLD[0].t10 259.254
R14879 WWLD[0] WWLD[0].n30 44.647
R14880 WWLD[0].n1 WWLD[0].n0 3.576
R14881 WWLD[0].n3 WWLD[0].n2 3.576
R14882 WWLD[0].n5 WWLD[0].n4 3.576
R14883 WWLD[0].n7 WWLD[0].n6 3.576
R14884 WWLD[0].n9 WWLD[0].n8 3.576
R14885 WWLD[0].n11 WWLD[0].n10 3.576
R14886 WWLD[0].n13 WWLD[0].n12 3.576
R14887 WWLD[0].n15 WWLD[0].n14 3.576
R14888 WWLD[0].n17 WWLD[0].n16 3.576
R14889 WWLD[0].n19 WWLD[0].n18 3.576
R14890 WWLD[0].n21 WWLD[0].n20 3.576
R14891 WWLD[0].n23 WWLD[0].n22 3.576
R14892 WWLD[0].n25 WWLD[0].n24 3.576
R14893 WWLD[0].n27 WWLD[0].n26 3.576
R14894 WWLD[0].n29 WWLD[0].n28 3.576
R14895 WWLD[0].n2 WWLD[0].n1 1.317
R14896 WWLD[0].n4 WWLD[0].n3 1.317
R14897 WWLD[0].n6 WWLD[0].n5 1.317
R14898 WWLD[0].n8 WWLD[0].n7 1.317
R14899 WWLD[0].n10 WWLD[0].n9 1.317
R14900 WWLD[0].n12 WWLD[0].n11 1.317
R14901 WWLD[0].n14 WWLD[0].n13 1.317
R14902 WWLD[0].n16 WWLD[0].n15 1.317
R14903 WWLD[0].n18 WWLD[0].n17 1.317
R14904 WWLD[0].n20 WWLD[0].n19 1.317
R14905 WWLD[0].n22 WWLD[0].n21 1.317
R14906 WWLD[0].n24 WWLD[0].n23 1.317
R14907 WWLD[0].n26 WWLD[0].n25 1.317
R14908 WWLD[0].n28 WWLD[0].n27 1.317
R14909 WWLD[0].n30 WWLD[0].n29 1.317
R14910 a_8902_4671.n0 a_8902_4671.t1 362.857
R14911 a_8902_4671.t4 a_8902_4671.t3 337.399
R14912 a_8902_4671.t3 a_8902_4671.t5 298.839
R14913 a_8902_4671.n0 a_8902_4671.t4 280.405
R14914 a_8902_4671.n1 a_8902_4671.t0 200
R14915 a_8902_4671.n1 a_8902_4671.n0 172.311
R14916 a_8902_4671.n2 a_8902_4671.n1 24
R14917 a_8902_4671.n1 a_8902_4671.t2 21.212
R14918 a_3152_3892.n0 a_3152_3892.t1 362.857
R14919 a_3152_3892.t4 a_3152_3892.t5 337.399
R14920 a_3152_3892.t5 a_3152_3892.t3 298.839
R14921 a_3152_3892.n0 a_3152_3892.t4 280.405
R14922 a_3152_3892.n1 a_3152_3892.t2 200
R14923 a_3152_3892.n1 a_3152_3892.n0 172.311
R14924 a_3152_3892.n2 a_3152_3892.n1 24
R14925 a_3152_3892.n1 a_3152_3892.t0 21.212
R14926 a_3165_3907.t0 a_3165_3907.t1 242.857
R14927 RWL[5].n0 RWL[5].t7 154.243
R14928 RWL[5].n14 RWL[5].t13 149.249
R14929 RWL[5].n13 RWL[5].t2 149.249
R14930 RWL[5].n12 RWL[5].t9 149.249
R14931 RWL[5].n11 RWL[5].t14 149.249
R14932 RWL[5].n10 RWL[5].t11 149.249
R14933 RWL[5].n9 RWL[5].t3 149.249
R14934 RWL[5].n8 RWL[5].t10 149.249
R14935 RWL[5].n7 RWL[5].t0 149.249
R14936 RWL[5].n6 RWL[5].t12 149.249
R14937 RWL[5].n5 RWL[5].t6 149.249
R14938 RWL[5].n4 RWL[5].t15 149.249
R14939 RWL[5].n3 RWL[5].t4 149.249
R14940 RWL[5].n2 RWL[5].t5 149.249
R14941 RWL[5].n1 RWL[5].t8 149.249
R14942 RWL[5].n0 RWL[5].t1 149.249
R14943 RWL[5] RWL[5].n14 42.872
R14944 RWL[5].n1 RWL[5].n0 4.994
R14945 RWL[5].n2 RWL[5].n1 4.994
R14946 RWL[5].n3 RWL[5].n2 4.994
R14947 RWL[5].n4 RWL[5].n3 4.994
R14948 RWL[5].n5 RWL[5].n4 4.994
R14949 RWL[5].n6 RWL[5].n5 4.994
R14950 RWL[5].n7 RWL[5].n6 4.994
R14951 RWL[5].n8 RWL[5].n7 4.994
R14952 RWL[5].n9 RWL[5].n8 4.994
R14953 RWL[5].n10 RWL[5].n9 4.994
R14954 RWL[5].n11 RWL[5].n10 4.994
R14955 RWL[5].n12 RWL[5].n11 4.994
R14956 RWL[5].n13 RWL[5].n12 4.994
R14957 RWL[5].n14 RWL[5].n13 4.994
R14958 a_4315_2421.t0 a_4315_2421.t1 242.857
R14959 a_11776_n7216.n0 a_11776_n7216.t3 1464.36
R14960 a_11776_n7216.n0 a_11776_n7216.t4 713.588
R14961 a_11776_n7216.n1 a_11776_n7216.t0 374.998
R14962 a_11776_n7216.n1 a_11776_n7216.t1 273.351
R14963 a_11776_n7216.n2 a_11776_n7216.n0 143.764
R14964 a_11776_n7216.t2 a_11776_n7216.n2 78.209
R14965 a_11776_n7216.n2 a_11776_n7216.n1 4.517
R14966 a_11549_n6503.n0 a_11549_n6503.t0 65.064
R14967 a_11549_n6503.n0 a_11549_n6503.t2 42.011
R14968 a_11549_n6503.t1 a_11549_n6503.n0 2.113
R14969 a_4448_n8026.n0 a_4448_n8026.t0 65.063
R14970 a_4448_n8026.n0 a_4448_n8026.t2 42.011
R14971 a_4448_n8026.t1 a_4448_n8026.n0 2.113
R14972 a_4302_678.n0 a_4302_678.t2 362.857
R14973 a_4302_678.t4 a_4302_678.t3 337.399
R14974 a_4302_678.t3 a_4302_678.t5 298.839
R14975 a_4302_678.n0 a_4302_678.t4 280.405
R14976 a_4302_678.n1 a_4302_678.t0 200
R14977 a_4302_678.n1 a_4302_678.n0 172.311
R14978 a_4302_678.n2 a_4302_678.n1 24
R14979 a_4302_678.n1 a_4302_678.t1 21.212
R14980 a_4397_693.n0 a_4397_693.t2 358.166
R14981 a_4397_693.t5 a_4397_693.t4 337.399
R14982 a_4397_693.t4 a_4397_693.t3 285.986
R14983 a_4397_693.n0 a_4397_693.t5 282.573
R14984 a_4397_693.n1 a_4397_693.t0 202.857
R14985 a_4397_693.n1 a_4397_693.n0 173.817
R14986 a_4397_693.n1 a_4397_693.t1 20.826
R14987 a_4397_693.n2 a_4397_693.n1 20.689
R14988 RWL[14].n0 RWL[14].t15 154.243
R14989 RWL[14].n14 RWL[14].t12 149.249
R14990 RWL[14].n13 RWL[14].t9 149.249
R14991 RWL[14].n12 RWL[14].t7 149.249
R14992 RWL[14].n11 RWL[14].t1 149.249
R14993 RWL[14].n10 RWL[14].t11 149.249
R14994 RWL[14].n9 RWL[14].t3 149.249
R14995 RWL[14].n8 RWL[14].t2 149.249
R14996 RWL[14].n7 RWL[14].t13 149.249
R14997 RWL[14].n6 RWL[14].t4 149.249
R14998 RWL[14].n5 RWL[14].t14 149.249
R14999 RWL[14].n4 RWL[14].t6 149.249
R15000 RWL[14].n3 RWL[14].t5 149.249
R15001 RWL[14].n2 RWL[14].t10 149.249
R15002 RWL[14].n1 RWL[14].t8 149.249
R15003 RWL[14].n0 RWL[14].t0 149.249
R15004 RWL[14] RWL[14].n14 42.872
R15005 RWL[14].n1 RWL[14].n0 4.994
R15006 RWL[14].n2 RWL[14].n1 4.994
R15007 RWL[14].n3 RWL[14].n2 4.994
R15008 RWL[14].n4 RWL[14].n3 4.994
R15009 RWL[14].n5 RWL[14].n4 4.994
R15010 RWL[14].n6 RWL[14].n5 4.994
R15011 RWL[14].n7 RWL[14].n6 4.994
R15012 RWL[14].n8 RWL[14].n7 4.994
R15013 RWL[14].n9 RWL[14].n8 4.994
R15014 RWL[14].n10 RWL[14].n9 4.994
R15015 RWL[14].n11 RWL[14].n10 4.994
R15016 RWL[14].n12 RWL[14].n11 4.994
R15017 RWL[14].n13 RWL[14].n12 4.994
R15018 RWL[14].n14 RWL[14].n13 4.994
R15019 a_8340_211.t0 a_8340_211.t1 242.857
R15020 a_5452_2928.n0 a_5452_2928.t1 362.857
R15021 a_5452_2928.t4 a_5452_2928.t5 337.399
R15022 a_5452_2928.t5 a_5452_2928.t3 298.839
R15023 a_5452_2928.n0 a_5452_2928.t4 280.405
R15024 a_5452_2928.n1 a_5452_2928.t2 200
R15025 a_5452_2928.n1 a_5452_2928.n0 172.311
R15026 a_5452_2928.n2 a_5452_2928.n1 24
R15027 a_5452_2928.n1 a_5452_2928.t0 21.212
R15028 a_5465_2943.t0 a_5465_2943.t1 242.857
R15029 a_7752_960.n0 a_7752_960.t1 362.857
R15030 a_7752_960.t3 a_7752_960.t5 337.399
R15031 a_7752_960.t5 a_7752_960.t4 298.839
R15032 a_7752_960.n0 a_7752_960.t3 280.405
R15033 a_7752_960.n1 a_7752_960.t0 200
R15034 a_7752_960.n1 a_7752_960.n0 172.311
R15035 a_7752_960.n2 a_7752_960.n1 24
R15036 a_7752_960.n1 a_7752_960.t2 21.212
R15037 a_7847_975.n0 a_7847_975.t2 358.166
R15038 a_7847_975.t4 a_7847_975.t5 337.399
R15039 a_7847_975.t5 a_7847_975.t3 285.986
R15040 a_7847_975.n0 a_7847_975.t4 282.573
R15041 a_7847_975.n1 a_7847_975.t0 202.857
R15042 a_7847_975.n1 a_7847_975.n0 173.817
R15043 a_7847_975.n1 a_7847_975.t1 20.826
R15044 a_7847_975.n2 a_7847_975.n1 20.689
R15045 a_2577_678.n0 a_2577_678.t1 362.857
R15046 a_2577_678.t4 a_2577_678.t3 337.399
R15047 a_2577_678.t3 a_2577_678.t5 298.839
R15048 a_2577_678.n0 a_2577_678.t4 280.405
R15049 a_2577_678.n1 a_2577_678.t2 200
R15050 a_2577_678.n1 a_2577_678.n0 172.311
R15051 a_2577_678.n2 a_2577_678.n1 24
R15052 a_2577_678.n1 a_2577_678.t0 21.212
R15053 a_n3495_n7203.n0 a_n3495_n7203.t0 63.08
R15054 a_n3495_n7203.t1 a_n3495_n7203.n0 41.306
R15055 a_n3495_n7203.n0 a_n3495_n7203.t2 2.251
R15056 a_n3357_n7203.t0 a_n3357_n7203.t1 68.741
R15057 a_7752_n286.n0 a_7752_n286.t2 362.857
R15058 a_7752_n286.t3 a_7752_n286.t4 337.399
R15059 a_7752_n286.t4 a_7752_n286.t5 298.839
R15060 a_7752_n286.n0 a_7752_n286.t3 280.405
R15061 a_7752_n286.n1 a_7752_n286.t0 200
R15062 a_7752_n286.n1 a_7752_n286.n0 172.311
R15063 a_7752_n286.n2 a_7752_n286.n1 24
R15064 a_7752_n286.n1 a_7752_n286.t1 21.212
R15065 a_10659_n4470.n0 a_10659_n4470.t0 63.08
R15066 a_10659_n4470.n0 a_10659_n4470.t2 41.305
R15067 a_10659_n4470.t1 a_10659_n4470.n0 2.251
R15068 a_10797_n4470.t0 a_10797_n4470.t1 68.741
R15069 a_4972_4686.n0 a_4972_4686.t2 358.166
R15070 a_4972_4686.t3 a_4972_4686.t5 337.399
R15071 a_4972_4686.t5 a_4972_4686.t4 285.986
R15072 a_4972_4686.n0 a_4972_4686.t3 282.573
R15073 a_4972_4686.n1 a_4972_4686.t0 202.857
R15074 a_4972_4686.n1 a_4972_4686.n0 173.817
R15075 a_4972_4686.n1 a_4972_4686.t1 20.826
R15076 a_4972_4686.n2 a_4972_4686.n1 20.689
R15077 a_4877_4671.n0 a_4877_4671.t1 362.857
R15078 a_4877_4671.t4 a_4877_4671.t3 337.399
R15079 a_4877_4671.t3 a_4877_4671.t5 298.839
R15080 a_4877_4671.n0 a_4877_4671.t4 280.405
R15081 a_4877_4671.n1 a_4877_4671.t2 200
R15082 a_4877_4671.n1 a_4877_4671.n0 172.311
R15083 a_4877_4671.n2 a_4877_4671.n1 24
R15084 a_4877_4671.n1 a_4877_4671.t0 21.212
R15085 a_3727_3410.n0 a_3727_3410.t2 362.857
R15086 a_3727_3410.t3 a_3727_3410.t4 337.399
R15087 a_3727_3410.t4 a_3727_3410.t5 298.839
R15088 a_3727_3410.n0 a_3727_3410.t3 280.405
R15089 a_3727_3410.n1 a_3727_3410.t0 200
R15090 a_3727_3410.n1 a_3727_3410.n0 172.311
R15091 a_3727_3410.n2 a_3727_3410.n1 24
R15092 a_3727_3410.n1 a_3727_3410.t1 21.212
R15093 a_3822_3425.n0 a_3822_3425.t2 358.166
R15094 a_3822_3425.t5 a_3822_3425.t4 337.399
R15095 a_3822_3425.t4 a_3822_3425.t3 285.986
R15096 a_3822_3425.n0 a_3822_3425.t5 282.573
R15097 a_3822_3425.n1 a_3822_3425.t0 202.857
R15098 a_3822_3425.n1 a_3822_3425.n0 173.817
R15099 a_3822_3425.n1 a_3822_3425.t1 20.826
R15100 a_3822_3425.n2 a_3822_3425.n1 20.689
R15101 a_7272_211.n0 a_7272_211.t0 358.166
R15102 a_7272_211.t4 a_7272_211.t3 337.399
R15103 a_7272_211.t3 a_7272_211.t5 285.986
R15104 a_7272_211.n0 a_7272_211.t4 282.573
R15105 a_7272_211.n1 a_7272_211.t1 202.857
R15106 a_7272_211.n1 a_7272_211.n0 173.817
R15107 a_7272_211.n1 a_7272_211.t2 20.826
R15108 a_7272_211.n2 a_7272_211.n1 20.689
R15109 a_7177_196.n0 a_7177_196.t2 362.857
R15110 a_7177_196.t4 a_7177_196.t3 337.399
R15111 a_7177_196.t3 a_7177_196.t5 298.839
R15112 a_7177_196.n0 a_7177_196.t4 280.405
R15113 a_7177_196.n1 a_7177_196.t0 200
R15114 a_7177_196.n1 a_7177_196.n0 172.311
R15115 a_7177_196.n2 a_7177_196.n1 24
R15116 a_7177_196.n1 a_7177_196.t1 21.212
R15117 a_1460_n1371.n1 a_1460_n1371.t3 550.94
R15118 a_1460_n1371.n1 a_1460_n1371.t4 500.621
R15119 a_1460_n1371.t2 a_1460_n1371.n2 192.787
R15120 a_1460_n1371.n0 a_1460_n1371.t0 163.997
R15121 a_1460_n1371.n2 a_1460_n1371.n1 149.035
R15122 a_1460_n1371.n0 a_1460_n1371.t1 54.068
R15123 a_1460_n1371.n2 a_1460_n1371.n0 17.317
R15124 a_1703_n1770.n0 a_1703_n1770.t1 160.619
R15125 a_1703_n1770.t0 a_1703_n1770.n0 151.153
R15126 SA_OUT[2].n1 SA_OUT[2].t3 661.027
R15127 SA_OUT[2].n1 SA_OUT[2].t4 392.255
R15128 SA_OUT[2].n2 SA_OUT[2].t1 223.716
R15129 SA_OUT[2].n0 SA_OUT[2].t0 153.977
R15130 SA_OUT[2].n2 SA_OUT[2].n1 143.764
R15131 SA_OUT[2].n0 SA_OUT[2].t2 59.86
R15132 SA_OUT[2] SA_OUT[2].n3 23.125
R15133 SA_OUT[2].n3 SA_OUT[2].n0 3.764
R15134 SA_OUT[2].n3 SA_OUT[2].n2 0.752
R15135 a_6492_2180.t0 a_6492_2180.t1 242.857
R15136 a_372_n271.n0 a_372_n271.t1 358.166
R15137 a_372_n271.t3 a_372_n271.t5 337.399
R15138 a_372_n271.t5 a_372_n271.t4 285.986
R15139 a_372_n271.n0 a_372_n271.t3 282.573
R15140 a_372_n271.n1 a_372_n271.t0 202.857
R15141 a_372_n271.n1 a_372_n271.n0 173.817
R15142 a_372_n271.n1 a_372_n271.t2 20.826
R15143 a_372_n271.n2 a_372_n271.n1 20.689
R15144 a_277_n286.n0 a_277_n286.t1 362.857
R15145 a_277_n286.t5 a_277_n286.t3 337.399
R15146 a_277_n286.t3 a_277_n286.t4 298.839
R15147 a_277_n286.n0 a_277_n286.t5 280.405
R15148 a_277_n286.n1 a_277_n286.t2 200
R15149 a_277_n286.n1 a_277_n286.n0 172.311
R15150 a_277_n286.n2 a_277_n286.n1 24
R15151 a_277_n286.n1 a_277_n286.t0 21.212
R15152 ADC13_OUT[0].n0 ADC13_OUT[0].t4 1354.27
R15153 ADC13_OUT[0].n0 ADC13_OUT[0].t3 821.954
R15154 ADC13_OUT[0].n3 ADC13_OUT[0].t0 328.315
R15155 ADC13_OUT[0].n2 ADC13_OUT[0].t1 266.575
R15156 ADC13_OUT[0].n1 ADC13_OUT[0].n0 149.035
R15157 ADC13_OUT[0] ADC13_OUT[0].n3 61.946
R15158 ADC13_OUT[0].n3 ADC13_OUT[0].n2 55.717
R15159 ADC13_OUT[0].n1 ADC13_OUT[0].t2 46.723
R15160 ADC13_OUT[0].n2 ADC13_OUT[0].n1 17.317
R15161 a_11776_n4483.n0 a_11776_n4483.t3 1464.36
R15162 a_11776_n4483.n0 a_11776_n4483.t4 713.588
R15163 a_11776_n4483.n1 a_11776_n4483.t0 374.998
R15164 a_11776_n4483.n1 a_11776_n4483.t1 273.351
R15165 a_11776_n4483.n2 a_11776_n4483.n0 143.764
R15166 a_11776_n4483.t2 a_11776_n4483.n2 78.209
R15167 a_11776_n4483.n2 a_11776_n4483.n1 4.517
R15168 Din[1].n0 Din[1].t0 215.292
R15169 Din[1].n0 Din[1].t1 187.376
R15170 Din[1] Din[1].n0 84.894
R15171 a_927_n2234.n2 a_927_n2234.t1 282.97
R15172 a_927_n2234.n1 a_927_n2234.t3 240.683
R15173 a_927_n2234.n0 a_927_n2234.t4 209.208
R15174 a_927_n2234.n0 a_927_n2234.t2 194.167
R15175 a_927_n2234.t0 a_927_n2234.n2 183.404
R15176 a_927_n2234.n1 a_927_n2234.n0 14.805
R15177 a_927_n2234.n2 a_927_n2234.n1 6.415
R15178 a_4890_n953.t42 a_4890_n953.n46 176.385
R15179 a_4890_n953.n22 a_4890_n953.t12 67.378
R15180 a_4890_n953.n0 a_4890_n953.t7 66.92
R15181 a_4890_n953.n1 a_4890_n953.t3 66.92
R15182 a_4890_n953.n2 a_4890_n953.t10 66.92
R15183 a_4890_n953.n3 a_4890_n953.t5 66.92
R15184 a_4890_n953.n4 a_4890_n953.t0 66.92
R15185 a_4890_n953.n5 a_4890_n953.t24 66.92
R15186 a_4890_n953.n6 a_4890_n953.t47 66.92
R15187 a_4890_n953.n7 a_4890_n953.t31 66.92
R15188 a_4890_n953.n8 a_4890_n953.t26 66.92
R15189 a_4890_n953.n9 a_4890_n953.t35 66.92
R15190 a_4890_n953.n10 a_4890_n953.t18 66.92
R15191 a_4890_n953.n11 a_4890_n953.t37 66.92
R15192 a_4890_n953.n12 a_4890_n953.t32 66.92
R15193 a_4890_n953.n13 a_4890_n953.t38 66.92
R15194 a_4890_n953.n14 a_4890_n953.t34 66.92
R15195 a_4890_n953.n15 a_4890_n953.t27 66.92
R15196 a_4890_n953.n16 a_4890_n953.t17 66.92
R15197 a_4890_n953.n17 a_4890_n953.t29 66.92
R15198 a_4890_n953.n18 a_4890_n953.t21 66.92
R15199 a_4890_n953.n19 a_4890_n953.t30 66.92
R15200 a_4890_n953.n20 a_4890_n953.t11 66.92
R15201 a_4890_n953.n21 a_4890_n953.t4 66.92
R15202 a_4890_n953.n22 a_4890_n953.t2 66.92
R15203 a_4890_n953.n23 a_4890_n953.t15 65.518
R15204 a_4890_n953.n45 a_4890_n953.t6 63.519
R15205 a_4890_n953.n44 a_4890_n953.t1 63.519
R15206 a_4890_n953.n43 a_4890_n953.t8 63.519
R15207 a_4890_n953.n42 a_4890_n953.t14 63.519
R15208 a_4890_n953.n41 a_4890_n953.t43 63.519
R15209 a_4890_n953.n40 a_4890_n953.t46 63.519
R15210 a_4890_n953.n39 a_4890_n953.t20 63.519
R15211 a_4890_n953.n38 a_4890_n953.t19 63.519
R15212 a_4890_n953.n37 a_4890_n953.t23 63.519
R15213 a_4890_n953.n36 a_4890_n953.t45 63.519
R15214 a_4890_n953.n35 a_4890_n953.t36 63.519
R15215 a_4890_n953.n34 a_4890_n953.t39 63.519
R15216 a_4890_n953.n33 a_4890_n953.t40 63.519
R15217 a_4890_n953.n32 a_4890_n953.t25 63.519
R15218 a_4890_n953.n31 a_4890_n953.t22 63.519
R15219 a_4890_n953.n30 a_4890_n953.t44 63.519
R15220 a_4890_n953.n29 a_4890_n953.t41 63.519
R15221 a_4890_n953.n28 a_4890_n953.t48 63.519
R15222 a_4890_n953.n27 a_4890_n953.t33 63.519
R15223 a_4890_n953.n26 a_4890_n953.t28 63.519
R15224 a_4890_n953.n25 a_4890_n953.t9 63.519
R15225 a_4890_n953.n24 a_4890_n953.t16 63.519
R15226 a_4890_n953.n23 a_4890_n953.t13 63.519
R15227 a_4890_n953.n46 a_4890_n953.n0 19.599
R15228 a_4890_n953.n46 a_4890_n953.n45 15.67
R15229 a_4890_n953.n44 a_4890_n953.n43 2.524
R15230 a_4890_n953.n24 a_4890_n953.n23 2.498
R15231 a_4890_n953.n21 a_4890_n953.n22 2.495
R15232 a_4890_n953.n1 a_4890_n953.n2 2.459
R15233 a_4890_n953.n38 a_4890_n953.n37 2.364
R15234 a_4890_n953.n30 a_4890_n953.n29 2.355
R15235 a_4890_n953.n7 a_4890_n953.n8 2.299
R15236 a_4890_n953.n15 a_4890_n953.n16 2.29
R15237 a_4890_n953.n16 a_4890_n953.n17 2.057
R15238 a_4890_n953.n8 a_4890_n953.n9 2.057
R15239 a_4890_n953.n2 a_4890_n953.n3 2.057
R15240 a_4890_n953.n0 a_4890_n953.n1 2.057
R15241 a_4890_n953.n45 a_4890_n953.n44 1.998
R15242 a_4890_n953.n43 a_4890_n953.n42 1.998
R15243 a_4890_n953.n42 a_4890_n953.n41 1.998
R15244 a_4890_n953.n41 a_4890_n953.n40 1.998
R15245 a_4890_n953.n40 a_4890_n953.n39 1.998
R15246 a_4890_n953.n39 a_4890_n953.n38 1.998
R15247 a_4890_n953.n37 a_4890_n953.n36 1.998
R15248 a_4890_n953.n36 a_4890_n953.n35 1.998
R15249 a_4890_n953.n35 a_4890_n953.n34 1.998
R15250 a_4890_n953.n34 a_4890_n953.n33 1.998
R15251 a_4890_n953.n33 a_4890_n953.n32 1.998
R15252 a_4890_n953.n32 a_4890_n953.n31 1.998
R15253 a_4890_n953.n31 a_4890_n953.n30 1.998
R15254 a_4890_n953.n29 a_4890_n953.n28 1.998
R15255 a_4890_n953.n28 a_4890_n953.n27 1.998
R15256 a_4890_n953.n27 a_4890_n953.n26 1.998
R15257 a_4890_n953.n26 a_4890_n953.n25 1.998
R15258 a_4890_n953.n25 a_4890_n953.n24 1.998
R15259 a_4890_n953.n20 a_4890_n953.n21 1.995
R15260 a_4890_n953.n19 a_4890_n953.n20 1.995
R15261 a_4890_n953.n18 a_4890_n953.n19 1.995
R15262 a_4890_n953.n17 a_4890_n953.n18 1.995
R15263 a_4890_n953.n14 a_4890_n953.n15 1.995
R15264 a_4890_n953.n13 a_4890_n953.n14 1.995
R15265 a_4890_n953.n12 a_4890_n953.n13 1.995
R15266 a_4890_n953.n11 a_4890_n953.n12 1.995
R15267 a_4890_n953.n10 a_4890_n953.n11 1.995
R15268 a_4890_n953.n9 a_4890_n953.n10 1.995
R15269 a_4890_n953.n6 a_4890_n953.n7 1.995
R15270 a_4890_n953.n5 a_4890_n953.n6 1.995
R15271 a_4890_n953.n4 a_4890_n953.n5 1.995
R15272 a_4890_n953.n3 a_4890_n953.n4 1.995
R15273 a_5342_4148.t0 a_5342_4148.t1 242.857
R15274 ADC2_OUT[2].n0 ADC2_OUT[2].t3 1354.27
R15275 ADC2_OUT[2].n0 ADC2_OUT[2].t4 821.954
R15276 ADC2_OUT[2].n3 ADC2_OUT[2].t0 347.138
R15277 ADC2_OUT[2].n2 ADC2_OUT[2].t1 266.575
R15278 ADC2_OUT[2].n1 ADC2_OUT[2].n0 149.035
R15279 ADC2_OUT[2].n1 ADC2_OUT[2].t2 46.723
R15280 ADC2_OUT[2] ADC2_OUT[2].n3 37.69
R15281 ADC2_OUT[2].n3 ADC2_OUT[2].n2 36.894
R15282 ADC2_OUT[2].n2 ADC2_OUT[2].n1 17.317
R15283 a_n1163_n7203.n0 a_n1163_n7203.t0 63.08
R15284 a_n1163_n7203.n0 a_n1163_n7203.t2 41.305
R15285 a_n1163_n7203.t1 a_n1163_n7203.n0 2.251
R15286 a_n1233_n7216.n0 a_n1233_n7216.t4 1464.36
R15287 a_n1233_n7216.n0 a_n1233_n7216.t3 713.588
R15288 a_n1233_n7216.n1 a_n1233_n7216.t0 374.998
R15289 a_n1233_n7216.n1 a_n1233_n7216.t1 273.351
R15290 a_n1233_n7216.n2 a_n1233_n7216.n0 143.764
R15291 a_n1233_n7216.t2 a_n1233_n7216.n2 78.209
R15292 a_n1233_n7216.n2 a_n1233_n7216.n1 4.517
R15293 a_8997_4686.n0 a_8997_4686.t2 358.166
R15294 a_8997_4686.t4 a_8997_4686.t5 337.399
R15295 a_8997_4686.t5 a_8997_4686.t3 285.986
R15296 a_8997_4686.n0 a_8997_4686.t4 282.573
R15297 a_8997_4686.n1 a_8997_4686.t0 202.857
R15298 a_8997_4686.n1 a_8997_4686.n0 173.817
R15299 a_8997_4686.n1 a_8997_4686.t1 20.826
R15300 a_8997_4686.n2 a_8997_4686.n1 20.689
R15301 a_9367_4686.t0 a_9367_4686.t1 242.857
R15302 a_5720_4887.n25 a_5720_4887.t27 561.971
R15303 a_5720_4887.n0 a_5720_4887.t26 449.944
R15304 a_5720_4887.t10 a_5720_4887.n25 108.636
R15305 a_5720_4887.n0 a_5720_4887.t25 74.821
R15306 a_5720_4887.n24 a_5720_4887.t17 63.519
R15307 a_5720_4887.n23 a_5720_4887.t15 63.519
R15308 a_5720_4887.n22 a_5720_4887.t4 63.519
R15309 a_5720_4887.n21 a_5720_4887.t11 63.519
R15310 a_5720_4887.n20 a_5720_4887.t20 63.519
R15311 a_5720_4887.n19 a_5720_4887.t13 63.519
R15312 a_5720_4887.n18 a_5720_4887.t14 63.519
R15313 a_5720_4887.n17 a_5720_4887.t8 63.519
R15314 a_5720_4887.n16 a_5720_4887.t3 63.519
R15315 a_5720_4887.n15 a_5720_4887.t6 63.519
R15316 a_5720_4887.n14 a_5720_4887.t18 63.519
R15317 a_5720_4887.n13 a_5720_4887.t0 63.519
R15318 a_5720_4887.n12 a_5720_4887.t12 63.519
R15319 a_5720_4887.n11 a_5720_4887.t23 63.519
R15320 a_5720_4887.n10 a_5720_4887.t9 63.519
R15321 a_5720_4887.n9 a_5720_4887.t19 63.519
R15322 a_5720_4887.n8 a_5720_4887.t16 63.519
R15323 a_5720_4887.n7 a_5720_4887.t2 63.519
R15324 a_5720_4887.n6 a_5720_4887.t1 63.519
R15325 a_5720_4887.n5 a_5720_4887.t24 63.519
R15326 a_5720_4887.n4 a_5720_4887.t7 63.519
R15327 a_5720_4887.n3 a_5720_4887.t21 63.519
R15328 a_5720_4887.n2 a_5720_4887.t22 63.519
R15329 a_5720_4887.n1 a_5720_4887.t5 63.519
R15330 a_5720_4887.n1 a_5720_4887.n0 8.619
R15331 a_5720_4887.n25 a_5720_4887.n24 2.946
R15332 a_5720_4887.n23 a_5720_4887.n22 2.524
R15333 a_5720_4887.n3 a_5720_4887.n2 2.498
R15334 a_5720_4887.n17 a_5720_4887.n16 2.364
R15335 a_5720_4887.n9 a_5720_4887.n8 2.355
R15336 a_5720_4887.n24 a_5720_4887.n23 1.998
R15337 a_5720_4887.n22 a_5720_4887.n21 1.998
R15338 a_5720_4887.n21 a_5720_4887.n20 1.998
R15339 a_5720_4887.n20 a_5720_4887.n19 1.998
R15340 a_5720_4887.n19 a_5720_4887.n18 1.998
R15341 a_5720_4887.n18 a_5720_4887.n17 1.998
R15342 a_5720_4887.n16 a_5720_4887.n15 1.998
R15343 a_5720_4887.n15 a_5720_4887.n14 1.998
R15344 a_5720_4887.n14 a_5720_4887.n13 1.998
R15345 a_5720_4887.n13 a_5720_4887.n12 1.998
R15346 a_5720_4887.n12 a_5720_4887.n11 1.998
R15347 a_5720_4887.n11 a_5720_4887.n10 1.998
R15348 a_5720_4887.n10 a_5720_4887.n9 1.998
R15349 a_5720_4887.n8 a_5720_4887.n7 1.998
R15350 a_5720_4887.n7 a_5720_4887.n6 1.998
R15351 a_5720_4887.n6 a_5720_4887.n5 1.998
R15352 a_5720_4887.n5 a_5720_4887.n4 1.998
R15353 a_5720_4887.n4 a_5720_4887.n3 1.998
R15354 a_5720_4887.n2 a_5720_4887.n1 1.998
R15355 a_5452_3169.n0 a_5452_3169.t0 362.857
R15356 a_5452_3169.t3 a_5452_3169.t4 337.399
R15357 a_5452_3169.t4 a_5452_3169.t5 298.839
R15358 a_5452_3169.n0 a_5452_3169.t3 280.405
R15359 a_5452_3169.n1 a_5452_3169.t2 200
R15360 a_5452_3169.n1 a_5452_3169.n0 172.311
R15361 a_5452_3169.n2 a_5452_3169.n1 24
R15362 a_5452_3169.n1 a_5452_3169.t1 21.212
R15363 RWLB[2].n0 RWLB[2].t15 154.228
R15364 RWLB[2].n14 RWLB[2].t0 149.249
R15365 RWLB[2].n13 RWLB[2].t2 149.249
R15366 RWLB[2].n12 RWLB[2].t13 149.249
R15367 RWLB[2].n11 RWLB[2].t7 149.249
R15368 RWLB[2].n10 RWLB[2].t1 149.249
R15369 RWLB[2].n9 RWLB[2].t4 149.249
R15370 RWLB[2].n8 RWLB[2].t5 149.249
R15371 RWLB[2].n7 RWLB[2].t10 149.249
R15372 RWLB[2].n6 RWLB[2].t3 149.249
R15373 RWLB[2].n5 RWLB[2].t8 149.249
R15374 RWLB[2].n4 RWLB[2].t9 149.249
R15375 RWLB[2].n3 RWLB[2].t14 149.249
R15376 RWLB[2].n2 RWLB[2].t6 149.249
R15377 RWLB[2].n1 RWLB[2].t12 149.249
R15378 RWLB[2].n0 RWLB[2].t11 149.249
R15379 RWLB[2] RWLB[2].n14 47.816
R15380 RWLB[2].n1 RWLB[2].n0 4.979
R15381 RWLB[2].n2 RWLB[2].n1 4.979
R15382 RWLB[2].n3 RWLB[2].n2 4.979
R15383 RWLB[2].n4 RWLB[2].n3 4.979
R15384 RWLB[2].n5 RWLB[2].n4 4.979
R15385 RWLB[2].n6 RWLB[2].n5 4.979
R15386 RWLB[2].n7 RWLB[2].n6 4.979
R15387 RWLB[2].n8 RWLB[2].n7 4.979
R15388 RWLB[2].n9 RWLB[2].n8 4.979
R15389 RWLB[2].n10 RWLB[2].n9 4.979
R15390 RWLB[2].n11 RWLB[2].n10 4.979
R15391 RWLB[2].n12 RWLB[2].n11 4.979
R15392 RWLB[2].n13 RWLB[2].n12 4.979
R15393 RWLB[2].n14 RWLB[2].n13 4.979
R15394 a_742_3184.t0 a_742_3184.t1 242.857
R15395 a_947_2421.n0 a_947_2421.t2 358.166
R15396 a_947_2421.t5 a_947_2421.t3 337.399
R15397 a_947_2421.t3 a_947_2421.t4 285.986
R15398 a_947_2421.n0 a_947_2421.t5 282.573
R15399 a_947_2421.n1 a_947_2421.t0 202.857
R15400 a_947_2421.n1 a_947_2421.n0 173.817
R15401 a_947_2421.n1 a_947_2421.t1 20.826
R15402 a_947_2421.n2 a_947_2421.n1 20.689
R15403 a_852_2406.n0 a_852_2406.t2 362.857
R15404 a_852_2406.t3 a_852_2406.t4 337.399
R15405 a_852_2406.t4 a_852_2406.t5 298.839
R15406 a_852_2406.n0 a_852_2406.t3 280.405
R15407 a_852_2406.n1 a_852_2406.t0 200
R15408 a_852_2406.n1 a_852_2406.n0 172.311
R15409 a_852_2406.n2 a_852_2406.n1 24
R15410 a_852_2406.n1 a_852_2406.t1 21.212
R15411 RWL[6].n0 RWL[6].t15 154.243
R15412 RWL[6].n14 RWL[6].t5 149.249
R15413 RWL[6].n13 RWL[6].t10 149.249
R15414 RWL[6].n12 RWL[6].t1 149.249
R15415 RWL[6].n11 RWL[6].t6 149.249
R15416 RWL[6].n10 RWL[6].t3 149.249
R15417 RWL[6].n9 RWL[6].t11 149.249
R15418 RWL[6].n8 RWL[6].t2 149.249
R15419 RWL[6].n7 RWL[6].t8 149.249
R15420 RWL[6].n6 RWL[6].t4 149.249
R15421 RWL[6].n5 RWL[6].t14 149.249
R15422 RWL[6].n4 RWL[6].t7 149.249
R15423 RWL[6].n3 RWL[6].t12 149.249
R15424 RWL[6].n2 RWL[6].t13 149.249
R15425 RWL[6].n1 RWL[6].t0 149.249
R15426 RWL[6].n0 RWL[6].t9 149.249
R15427 RWL[6] RWL[6].n14 42.872
R15428 RWL[6].n1 RWL[6].n0 4.994
R15429 RWL[6].n2 RWL[6].n1 4.994
R15430 RWL[6].n3 RWL[6].n2 4.994
R15431 RWL[6].n4 RWL[6].n3 4.994
R15432 RWL[6].n5 RWL[6].n4 4.994
R15433 RWL[6].n6 RWL[6].n5 4.994
R15434 RWL[6].n7 RWL[6].n6 4.994
R15435 RWL[6].n8 RWL[6].n7 4.994
R15436 RWL[6].n9 RWL[6].n8 4.994
R15437 RWL[6].n10 RWL[6].n9 4.994
R15438 RWL[6].n11 RWL[6].n10 4.994
R15439 RWL[6].n12 RWL[6].n11 4.994
R15440 RWL[6].n13 RWL[6].n12 4.994
R15441 RWL[6].n14 RWL[6].n13 4.994
R15442 a_7765_2180.t0 a_7765_2180.t1 242.857
R15443 a_7765_n953.t46 a_7765_n953.n46 176.385
R15444 a_7765_n953.n22 a_7765_n953.t5 67.378
R15445 a_7765_n953.n0 a_7765_n953.t3 66.92
R15446 a_7765_n953.n1 a_7765_n953.t17 66.92
R15447 a_7765_n953.n2 a_7765_n953.t15 66.92
R15448 a_7765_n953.n3 a_7765_n953.t12 66.92
R15449 a_7765_n953.n4 a_7765_n953.t1 66.92
R15450 a_7765_n953.n5 a_7765_n953.t25 66.92
R15451 a_7765_n953.n6 a_7765_n953.t48 66.92
R15452 a_7765_n953.n7 a_7765_n953.t32 66.92
R15453 a_7765_n953.n8 a_7765_n953.t27 66.92
R15454 a_7765_n953.n9 a_7765_n953.t38 66.92
R15455 a_7765_n953.n10 a_7765_n953.t19 66.92
R15456 a_7765_n953.n11 a_7765_n953.t42 66.92
R15457 a_7765_n953.n12 a_7765_n953.t33 66.92
R15458 a_7765_n953.n13 a_7765_n953.t37 66.92
R15459 a_7765_n953.n14 a_7765_n953.t36 66.92
R15460 a_7765_n953.n15 a_7765_n953.t28 66.92
R15461 a_7765_n953.n16 a_7765_n953.t18 66.92
R15462 a_7765_n953.n17 a_7765_n953.t30 66.92
R15463 a_7765_n953.n18 a_7765_n953.t22 66.92
R15464 a_7765_n953.n19 a_7765_n953.t31 66.92
R15465 a_7765_n953.n20 a_7765_n953.t7 66.92
R15466 a_7765_n953.n21 a_7765_n953.t16 66.92
R15467 a_7765_n953.n22 a_7765_n953.t13 66.92
R15468 a_7765_n953.n23 a_7765_n953.t4 65.518
R15469 a_7765_n953.n45 a_7765_n953.t6 63.519
R15470 a_7765_n953.n44 a_7765_n953.t2 63.519
R15471 a_7765_n953.n43 a_7765_n953.t14 63.519
R15472 a_7765_n953.n42 a_7765_n953.t9 63.519
R15473 a_7765_n953.n41 a_7765_n953.t41 63.519
R15474 a_7765_n953.n40 a_7765_n953.t47 63.519
R15475 a_7765_n953.n39 a_7765_n953.t21 63.519
R15476 a_7765_n953.n38 a_7765_n953.t20 63.519
R15477 a_7765_n953.n37 a_7765_n953.t24 63.519
R15478 a_7765_n953.n36 a_7765_n953.t45 63.519
R15479 a_7765_n953.n35 a_7765_n953.t39 63.519
R15480 a_7765_n953.n34 a_7765_n953.t35 63.519
R15481 a_7765_n953.n33 a_7765_n953.t0 63.519
R15482 a_7765_n953.n32 a_7765_n953.t26 63.519
R15483 a_7765_n953.n31 a_7765_n953.t23 63.519
R15484 a_7765_n953.n30 a_7765_n953.t44 63.519
R15485 a_7765_n953.n29 a_7765_n953.t43 63.519
R15486 a_7765_n953.n28 a_7765_n953.t40 63.519
R15487 a_7765_n953.n27 a_7765_n953.t34 63.519
R15488 a_7765_n953.n26 a_7765_n953.t29 63.519
R15489 a_7765_n953.n25 a_7765_n953.t11 63.519
R15490 a_7765_n953.n24 a_7765_n953.t10 63.519
R15491 a_7765_n953.n23 a_7765_n953.t8 63.519
R15492 a_7765_n953.n46 a_7765_n953.n45 18.144
R15493 a_7765_n953.n46 a_7765_n953.n0 17.125
R15494 a_7765_n953.n44 a_7765_n953.n43 2.524
R15495 a_7765_n953.n24 a_7765_n953.n23 2.498
R15496 a_7765_n953.n21 a_7765_n953.n22 2.495
R15497 a_7765_n953.n1 a_7765_n953.n2 2.459
R15498 a_7765_n953.n38 a_7765_n953.n37 2.364
R15499 a_7765_n953.n30 a_7765_n953.n29 2.355
R15500 a_7765_n953.n7 a_7765_n953.n8 2.299
R15501 a_7765_n953.n15 a_7765_n953.n16 2.29
R15502 a_7765_n953.n16 a_7765_n953.n17 2.057
R15503 a_7765_n953.n8 a_7765_n953.n9 2.057
R15504 a_7765_n953.n2 a_7765_n953.n3 2.057
R15505 a_7765_n953.n0 a_7765_n953.n1 2.057
R15506 a_7765_n953.n45 a_7765_n953.n44 1.998
R15507 a_7765_n953.n43 a_7765_n953.n42 1.998
R15508 a_7765_n953.n42 a_7765_n953.n41 1.998
R15509 a_7765_n953.n41 a_7765_n953.n40 1.998
R15510 a_7765_n953.n40 a_7765_n953.n39 1.998
R15511 a_7765_n953.n39 a_7765_n953.n38 1.998
R15512 a_7765_n953.n37 a_7765_n953.n36 1.998
R15513 a_7765_n953.n36 a_7765_n953.n35 1.998
R15514 a_7765_n953.n35 a_7765_n953.n34 1.998
R15515 a_7765_n953.n34 a_7765_n953.n33 1.998
R15516 a_7765_n953.n33 a_7765_n953.n32 1.998
R15517 a_7765_n953.n32 a_7765_n953.n31 1.998
R15518 a_7765_n953.n31 a_7765_n953.n30 1.998
R15519 a_7765_n953.n29 a_7765_n953.n28 1.998
R15520 a_7765_n953.n28 a_7765_n953.n27 1.998
R15521 a_7765_n953.n27 a_7765_n953.n26 1.998
R15522 a_7765_n953.n26 a_7765_n953.n25 1.998
R15523 a_7765_n953.n25 a_7765_n953.n24 1.998
R15524 a_7765_n953.n20 a_7765_n953.n21 1.995
R15525 a_7765_n953.n19 a_7765_n953.n20 1.995
R15526 a_7765_n953.n18 a_7765_n953.n19 1.995
R15527 a_7765_n953.n17 a_7765_n953.n18 1.995
R15528 a_7765_n953.n14 a_7765_n953.n15 1.995
R15529 a_7765_n953.n13 a_7765_n953.n14 1.995
R15530 a_7765_n953.n12 a_7765_n953.n13 1.995
R15531 a_7765_n953.n11 a_7765_n953.n12 1.995
R15532 a_7765_n953.n10 a_7765_n953.n11 1.995
R15533 a_7765_n953.n9 a_7765_n953.n10 1.995
R15534 a_7765_n953.n6 a_7765_n953.n7 1.995
R15535 a_7765_n953.n5 a_7765_n953.n6 1.995
R15536 a_7765_n953.n4 a_7765_n953.n5 1.995
R15537 a_7765_n953.n3 a_7765_n953.n4 1.995
R15538 a_1502_n2234.n2 a_1502_n2234.t1 282.97
R15539 a_1502_n2234.n1 a_1502_n2234.t2 240.683
R15540 a_1502_n2234.n0 a_1502_n2234.t3 209.208
R15541 a_1502_n2234.n0 a_1502_n2234.t4 194.167
R15542 a_1502_n2234.t0 a_1502_n2234.n2 183.404
R15543 a_1502_n2234.n1 a_1502_n2234.n0 14.805
R15544 a_1502_n2234.n2 a_1502_n2234.n1 6.415
R15545 a_1743_n2086.t0 a_1743_n2086.t1 34.8
R15546 a_6615_4148.t0 a_6615_4148.t1 242.857
R15547 a_1522_2943.n0 a_1522_2943.t1 358.166
R15548 a_1522_2943.t5 a_1522_2943.t4 337.399
R15549 a_1522_2943.t4 a_1522_2943.t3 285.986
R15550 a_1522_2943.n0 a_1522_2943.t5 282.573
R15551 a_1522_2943.n1 a_1522_2943.t0 202.857
R15552 a_1522_2943.n1 a_1522_2943.n0 173.817
R15553 a_1522_2943.n1 a_1522_2943.t2 20.826
R15554 a_1522_2943.n2 a_1522_2943.n1 20.689
R15555 a_1892_2943.t0 a_1892_2943.t1 242.857
R15556 Iref0.n0 Iref0.t10 466.061
R15557 Iref0.n14 Iref0.t9 456.909
R15558 Iref0.n13 Iref0.t2 456.909
R15559 Iref0.n12 Iref0.t11 456.909
R15560 Iref0.n11 Iref0.t1 456.909
R15561 Iref0.n10 Iref0.t0 456.909
R15562 Iref0.n9 Iref0.t4 456.909
R15563 Iref0.n8 Iref0.t7 456.909
R15564 Iref0.n7 Iref0.t14 456.909
R15565 Iref0.n6 Iref0.t6 456.909
R15566 Iref0.n5 Iref0.t13 456.909
R15567 Iref0.n4 Iref0.t5 456.909
R15568 Iref0.n3 Iref0.t12 456.909
R15569 Iref0.n2 Iref0.t15 456.909
R15570 Iref0.n1 Iref0.t8 456.909
R15571 Iref0.n0 Iref0.t3 456.909
R15572 Iref0 Iref0.n14 39.584
R15573 Iref0.n12 Iref0.n11 8.671
R15574 Iref0.n13 Iref0.n12 8.671
R15575 Iref0.n10 Iref0.n9 8.649
R15576 Iref0.n11 Iref0.n10 8.649
R15577 Iref0.n1 Iref0.n0 8.634
R15578 Iref0.n4 Iref0.n3 8.634
R15579 Iref0.n5 Iref0.n4 8.634
R15580 Iref0.n6 Iref0.n5 8.634
R15581 Iref0.n7 Iref0.n6 8.634
R15582 Iref0.n8 Iref0.n7 8.634
R15583 Iref0.n9 Iref0.n8 8.634
R15584 Iref0.n2 Iref0.n1 8.627
R15585 Iref0.n3 Iref0.n2 8.627
R15586 Iref0.n14 Iref0.n13 6.561
R15587 a_9672_n4114.t1 a_9672_n4114.t0 336.812
R15588 a_372_3425.n0 a_372_3425.t1 358.166
R15589 a_372_3425.t3 a_372_3425.t5 337.399
R15590 a_372_3425.t5 a_372_3425.t4 285.986
R15591 a_372_3425.n0 a_372_3425.t3 282.573
R15592 a_372_3425.n1 a_372_3425.t0 202.857
R15593 a_372_3425.n1 a_372_3425.n0 173.817
R15594 a_372_3425.n1 a_372_3425.t2 20.826
R15595 a_372_3425.n2 a_372_3425.n1 20.689
R15596 a_277_3410.n0 a_277_3410.t1 362.857
R15597 a_277_3410.t3 a_277_3410.t4 337.399
R15598 a_277_3410.t4 a_277_3410.t5 298.839
R15599 a_277_3410.n0 a_277_3410.t3 280.405
R15600 a_277_3410.n1 a_277_3410.t2 200
R15601 a_277_3410.n1 a_277_3410.n0 172.311
R15602 a_277_3410.n2 a_277_3410.n1 24
R15603 a_277_3410.n1 a_277_3410.t0 21.212
R15604 a_2577_3651.n0 a_2577_3651.t1 362.857
R15605 a_2577_3651.t4 a_2577_3651.t5 337.399
R15606 a_2577_3651.t5 a_2577_3651.t3 298.839
R15607 a_2577_3651.n0 a_2577_3651.t4 280.405
R15608 a_2577_3651.n1 a_2577_3651.t2 200
R15609 a_2577_3651.n1 a_2577_3651.n0 172.311
R15610 a_2577_3651.n2 a_2577_3651.n1 24
R15611 a_2577_3651.n1 a_2577_3651.t0 21.212
R15612 a_2590_3666.t0 a_2590_3666.t1 242.857
R15613 a_n1233_n4483.n0 a_n1233_n4483.t4 1464.36
R15614 a_n1233_n4483.n0 a_n1233_n4483.t3 713.588
R15615 a_n1233_n4483.n1 a_n1233_n4483.t0 374.998
R15616 a_n1233_n4483.n1 a_n1233_n4483.t2 273.351
R15617 a_n1233_n4483.n2 a_n1233_n4483.n0 143.764
R15618 a_n1233_n4483.t1 a_n1233_n4483.n2 78.209
R15619 a_n1233_n4483.n2 a_n1233_n4483.n1 4.517
R15620 ADC2_OUT[0].n0 ADC2_OUT[0].t3 1354.27
R15621 ADC2_OUT[0].n0 ADC2_OUT[0].t4 821.954
R15622 ADC2_OUT[0].n3 ADC2_OUT[0].t0 344.126
R15623 ADC2_OUT[0].n2 ADC2_OUT[0].t1 266.575
R15624 ADC2_OUT[0].n1 ADC2_OUT[0].n0 149.035
R15625 ADC2_OUT[0] ADC2_OUT[0].n3 61.433
R15626 ADC2_OUT[0].n1 ADC2_OUT[0].t2 46.723
R15627 ADC2_OUT[0].n3 ADC2_OUT[0].n2 39.905
R15628 ADC2_OUT[0].n2 ADC2_OUT[0].n1 17.317
R15629 PRE_SRAM.n45 PRE_SRAM.t31 303.489
R15630 PRE_SRAM.n42 PRE_SRAM.t36 303.489
R15631 PRE_SRAM.n39 PRE_SRAM.t21 303.489
R15632 PRE_SRAM.n36 PRE_SRAM.t43 303.489
R15633 PRE_SRAM.n33 PRE_SRAM.t17 303.489
R15634 PRE_SRAM.n30 PRE_SRAM.t40 303.489
R15635 PRE_SRAM.n27 PRE_SRAM.t25 303.489
R15636 PRE_SRAM.n24 PRE_SRAM.t3 303.489
R15637 PRE_SRAM.n21 PRE_SRAM.t37 303.489
R15638 PRE_SRAM.n18 PRE_SRAM.t45 303.489
R15639 PRE_SRAM.n15 PRE_SRAM.t46 303.489
R15640 PRE_SRAM.n12 PRE_SRAM.t8 303.489
R15641 PRE_SRAM.n9 PRE_SRAM.t42 303.489
R15642 PRE_SRAM.n6 PRE_SRAM.t18 303.489
R15643 PRE_SRAM.n3 PRE_SRAM.t6 303.489
R15644 PRE_SRAM.n0 PRE_SRAM.t26 303.489
R15645 PRE_SRAM.n0 PRE_SRAM.t12 156.336
R15646 PRE_SRAM.n46 PRE_SRAM.t33 155.676
R15647 PRE_SRAM.n44 PRE_SRAM.t1 155.676
R15648 PRE_SRAM.n43 PRE_SRAM.t39 155.676
R15649 PRE_SRAM.n41 PRE_SRAM.t19 155.676
R15650 PRE_SRAM.n40 PRE_SRAM.t24 155.676
R15651 PRE_SRAM.n38 PRE_SRAM.t38 155.676
R15652 PRE_SRAM.n37 PRE_SRAM.t2 155.676
R15653 PRE_SRAM.n35 PRE_SRAM.t27 155.676
R15654 PRE_SRAM.n34 PRE_SRAM.t22 155.676
R15655 PRE_SRAM.n32 PRE_SRAM.t34 155.676
R15656 PRE_SRAM.n31 PRE_SRAM.t44 155.676
R15657 PRE_SRAM.n29 PRE_SRAM.t23 155.676
R15658 PRE_SRAM.n28 PRE_SRAM.t29 155.676
R15659 PRE_SRAM.n26 PRE_SRAM.t14 155.676
R15660 PRE_SRAM.n25 PRE_SRAM.t7 155.676
R15661 PRE_SRAM.n23 PRE_SRAM.t32 155.676
R15662 PRE_SRAM.n22 PRE_SRAM.t41 155.676
R15663 PRE_SRAM.n20 PRE_SRAM.t11 155.676
R15664 PRE_SRAM.n19 PRE_SRAM.t4 155.676
R15665 PRE_SRAM.n17 PRE_SRAM.t28 155.676
R15666 PRE_SRAM.n16 PRE_SRAM.t5 155.676
R15667 PRE_SRAM.n14 PRE_SRAM.t16 155.676
R15668 PRE_SRAM.n13 PRE_SRAM.t13 155.676
R15669 PRE_SRAM.n11 PRE_SRAM.t35 155.676
R15670 PRE_SRAM.n10 PRE_SRAM.t47 155.676
R15671 PRE_SRAM.n8 PRE_SRAM.t15 155.676
R15672 PRE_SRAM.n7 PRE_SRAM.t9 155.676
R15673 PRE_SRAM.n5 PRE_SRAM.t0 155.676
R15674 PRE_SRAM.n4 PRE_SRAM.t10 155.676
R15675 PRE_SRAM.n2 PRE_SRAM.t20 155.676
R15676 PRE_SRAM.n1 PRE_SRAM.t30 155.676
R15677 PRE_SRAM PRE_SRAM.n46 44.577
R15678 PRE_SRAM.n2 PRE_SRAM.n1 3.463
R15679 PRE_SRAM.n5 PRE_SRAM.n4 3.463
R15680 PRE_SRAM.n8 PRE_SRAM.n7 3.463
R15681 PRE_SRAM.n11 PRE_SRAM.n10 3.463
R15682 PRE_SRAM.n14 PRE_SRAM.n13 3.463
R15683 PRE_SRAM.n17 PRE_SRAM.n16 3.463
R15684 PRE_SRAM.n20 PRE_SRAM.n19 3.463
R15685 PRE_SRAM.n23 PRE_SRAM.n22 3.463
R15686 PRE_SRAM.n26 PRE_SRAM.n25 3.463
R15687 PRE_SRAM.n29 PRE_SRAM.n28 3.463
R15688 PRE_SRAM.n32 PRE_SRAM.n31 3.463
R15689 PRE_SRAM.n35 PRE_SRAM.n34 3.463
R15690 PRE_SRAM.n38 PRE_SRAM.n37 3.463
R15691 PRE_SRAM.n41 PRE_SRAM.n40 3.463
R15692 PRE_SRAM.n44 PRE_SRAM.n43 3.463
R15693 PRE_SRAM.n1 PRE_SRAM.n0 0.66
R15694 PRE_SRAM.n3 PRE_SRAM.n2 0.66
R15695 PRE_SRAM.n4 PRE_SRAM.n3 0.66
R15696 PRE_SRAM.n6 PRE_SRAM.n5 0.66
R15697 PRE_SRAM.n7 PRE_SRAM.n6 0.66
R15698 PRE_SRAM.n9 PRE_SRAM.n8 0.66
R15699 PRE_SRAM.n10 PRE_SRAM.n9 0.66
R15700 PRE_SRAM.n12 PRE_SRAM.n11 0.66
R15701 PRE_SRAM.n13 PRE_SRAM.n12 0.66
R15702 PRE_SRAM.n15 PRE_SRAM.n14 0.66
R15703 PRE_SRAM.n16 PRE_SRAM.n15 0.66
R15704 PRE_SRAM.n18 PRE_SRAM.n17 0.66
R15705 PRE_SRAM.n19 PRE_SRAM.n18 0.66
R15706 PRE_SRAM.n21 PRE_SRAM.n20 0.66
R15707 PRE_SRAM.n22 PRE_SRAM.n21 0.66
R15708 PRE_SRAM.n24 PRE_SRAM.n23 0.66
R15709 PRE_SRAM.n25 PRE_SRAM.n24 0.66
R15710 PRE_SRAM.n27 PRE_SRAM.n26 0.66
R15711 PRE_SRAM.n28 PRE_SRAM.n27 0.66
R15712 PRE_SRAM.n30 PRE_SRAM.n29 0.66
R15713 PRE_SRAM.n31 PRE_SRAM.n30 0.66
R15714 PRE_SRAM.n33 PRE_SRAM.n32 0.66
R15715 PRE_SRAM.n34 PRE_SRAM.n33 0.66
R15716 PRE_SRAM.n36 PRE_SRAM.n35 0.66
R15717 PRE_SRAM.n37 PRE_SRAM.n36 0.66
R15718 PRE_SRAM.n39 PRE_SRAM.n38 0.66
R15719 PRE_SRAM.n40 PRE_SRAM.n39 0.66
R15720 PRE_SRAM.n42 PRE_SRAM.n41 0.66
R15721 PRE_SRAM.n43 PRE_SRAM.n42 0.66
R15722 PRE_SRAM.n45 PRE_SRAM.n44 0.66
R15723 PRE_SRAM.n46 PRE_SRAM.n45 0.66
R15724 a_4877_3651.n0 a_4877_3651.t1 362.857
R15725 a_4877_3651.t3 a_4877_3651.t5 337.399
R15726 a_4877_3651.t5 a_4877_3651.t4 298.839
R15727 a_4877_3651.n0 a_4877_3651.t3 280.405
R15728 a_4877_3651.n1 a_4877_3651.t2 200
R15729 a_4877_3651.n1 a_4877_3651.n0 172.311
R15730 a_4877_3651.n2 a_4877_3651.n1 24
R15731 a_4877_3651.n1 a_4877_3651.t0 21.212
R15732 a_4972_3666.n0 a_4972_3666.t1 358.166
R15733 a_4972_3666.t4 a_4972_3666.t3 337.399
R15734 a_4972_3666.t3 a_4972_3666.t5 285.986
R15735 a_4972_3666.n0 a_4972_3666.t4 282.573
R15736 a_4972_3666.n1 a_4972_3666.t2 202.857
R15737 a_4972_3666.n1 a_4972_3666.n0 173.817
R15738 a_4972_3666.n1 a_4972_3666.t0 20.826
R15739 a_4972_3666.n2 a_4972_3666.n1 20.689
R15740 a_2002_1201.n0 a_2002_1201.t0 362.857
R15741 a_2002_1201.t3 a_2002_1201.t5 337.399
R15742 a_2002_1201.t5 a_2002_1201.t4 298.839
R15743 a_2002_1201.n0 a_2002_1201.t3 280.405
R15744 a_2002_1201.n1 a_2002_1201.t2 200
R15745 a_2002_1201.n1 a_2002_1201.n0 172.311
R15746 a_2002_1201.n2 a_2002_1201.n1 24
R15747 a_2002_1201.n1 a_2002_1201.t1 21.212
R15748 a_2097_1216.n0 a_2097_1216.t2 358.166
R15749 a_2097_1216.t5 a_2097_1216.t3 337.399
R15750 a_2097_1216.t3 a_2097_1216.t4 285.986
R15751 a_2097_1216.n0 a_2097_1216.t5 282.573
R15752 a_2097_1216.n1 a_2097_1216.t0 202.857
R15753 a_2097_1216.n1 a_2097_1216.n0 173.817
R15754 a_2097_1216.n1 a_2097_1216.t1 20.826
R15755 a_2097_1216.n2 a_2097_1216.n1 20.689
R15756 a_7847_452.n0 a_7847_452.t2 358.166
R15757 a_7847_452.t3 a_7847_452.t5 337.399
R15758 a_7847_452.t5 a_7847_452.t4 285.986
R15759 a_7847_452.n0 a_7847_452.t3 282.573
R15760 a_7847_452.n1 a_7847_452.t0 202.857
R15761 a_7847_452.n1 a_7847_452.n0 173.817
R15762 a_7847_452.n1 a_7847_452.t1 20.826
R15763 a_7847_452.n2 a_7847_452.n1 20.689
R15764 a_8217_n812.t0 a_8217_n812.t1 242.857
R15765 a_1892_975.t0 a_1892_975.t1 242.857
R15766 a_8433_n953.n25 a_8433_n953.t27 561.971
R15767 a_8433_n953.n0 a_8433_n953.t4 461.908
R15768 a_8433_n953.t12 a_8433_n953.n25 108.635
R15769 a_8433_n953.n0 a_8433_n953.t3 79.512
R15770 a_8433_n953.n24 a_8433_n953.t19 65.401
R15771 a_8433_n953.n23 a_8433_n953.t17 65.401
R15772 a_8433_n953.n22 a_8433_n953.t7 65.401
R15773 a_8433_n953.n21 a_8433_n953.t13 65.401
R15774 a_8433_n953.n20 a_8433_n953.t22 65.401
R15775 a_8433_n953.n19 a_8433_n953.t15 65.401
R15776 a_8433_n953.n18 a_8433_n953.t16 65.401
R15777 a_8433_n953.n17 a_8433_n953.t11 65.401
R15778 a_8433_n953.n16 a_8433_n953.t2 65.401
R15779 a_8433_n953.n15 a_8433_n953.t9 65.401
R15780 a_8433_n953.n14 a_8433_n953.t20 65.401
R15781 a_8433_n953.n13 a_8433_n953.t5 65.401
R15782 a_8433_n953.n12 a_8433_n953.t14 65.401
R15783 a_8433_n953.n11 a_8433_n953.t25 65.401
R15784 a_8433_n953.n10 a_8433_n953.t6 65.401
R15785 a_8433_n953.n9 a_8433_n953.t21 65.401
R15786 a_8433_n953.n8 a_8433_n953.t18 65.401
R15787 a_8433_n953.n7 a_8433_n953.t1 65.401
R15788 a_8433_n953.n6 a_8433_n953.t0 65.401
R15789 a_8433_n953.n5 a_8433_n953.t26 65.401
R15790 a_8433_n953.n4 a_8433_n953.t10 65.401
R15791 a_8433_n953.n3 a_8433_n953.t23 65.401
R15792 a_8433_n953.n2 a_8433_n953.t24 65.401
R15793 a_8433_n953.n1 a_8433_n953.t8 65.401
R15794 a_8433_n953.n1 a_8433_n953.n0 5.64
R15795 a_8433_n953.n25 a_8433_n953.n24 4.438
R15796 a_8433_n953.n23 a_8433_n953.n22 2.524
R15797 a_8433_n953.n3 a_8433_n953.n2 2.498
R15798 a_8433_n953.n17 a_8433_n953.n16 2.364
R15799 a_8433_n953.n9 a_8433_n953.n8 2.355
R15800 a_8433_n953.n2 a_8433_n953.n1 1.998
R15801 a_8433_n953.n4 a_8433_n953.n3 1.998
R15802 a_8433_n953.n5 a_8433_n953.n4 1.998
R15803 a_8433_n953.n6 a_8433_n953.n5 1.998
R15804 a_8433_n953.n7 a_8433_n953.n6 1.998
R15805 a_8433_n953.n8 a_8433_n953.n7 1.998
R15806 a_8433_n953.n10 a_8433_n953.n9 1.998
R15807 a_8433_n953.n11 a_8433_n953.n10 1.998
R15808 a_8433_n953.n12 a_8433_n953.n11 1.998
R15809 a_8433_n953.n13 a_8433_n953.n12 1.998
R15810 a_8433_n953.n14 a_8433_n953.n13 1.998
R15811 a_8433_n953.n15 a_8433_n953.n14 1.998
R15812 a_8433_n953.n16 a_8433_n953.n15 1.998
R15813 a_8433_n953.n18 a_8433_n953.n17 1.998
R15814 a_8433_n953.n19 a_8433_n953.n18 1.998
R15815 a_8433_n953.n20 a_8433_n953.n19 1.998
R15816 a_8433_n953.n21 a_8433_n953.n20 1.998
R15817 a_8433_n953.n22 a_8433_n953.n21 1.998
R15818 a_8433_n953.n24 a_8433_n953.n23 1.998
R15819 a_5547_3184.n0 a_5547_3184.t2 358.166
R15820 a_5547_3184.t4 a_5547_3184.t5 337.399
R15821 a_5547_3184.t5 a_5547_3184.t3 285.986
R15822 a_5547_3184.n0 a_5547_3184.t4 282.573
R15823 a_5547_3184.n1 a_5547_3184.t0 202.857
R15824 a_5547_3184.n1 a_5547_3184.n0 173.817
R15825 a_5547_3184.n1 a_5547_3184.t1 20.826
R15826 a_5547_3184.n2 a_5547_3184.n1 20.689
R15827 a_5917_3184.t0 a_5917_3184.t1 242.857
R15828 a_7272_3425.n0 a_7272_3425.t1 358.166
R15829 a_7272_3425.t3 a_7272_3425.t5 337.399
R15830 a_7272_3425.t5 a_7272_3425.t4 285.986
R15831 a_7272_3425.n0 a_7272_3425.t3 282.573
R15832 a_7272_3425.n1 a_7272_3425.t0 202.857
R15833 a_7272_3425.n1 a_7272_3425.n0 173.817
R15834 a_7272_3425.n1 a_7272_3425.t2 20.826
R15835 a_7272_3425.n2 a_7272_3425.n1 20.689
R15836 a_6602_3892.n0 a_6602_3892.t1 362.857
R15837 a_6602_3892.t5 a_6602_3892.t4 337.399
R15838 a_6602_3892.t4 a_6602_3892.t3 298.839
R15839 a_6602_3892.n0 a_6602_3892.t5 280.405
R15840 a_6602_3892.n1 a_6602_3892.t2 200
R15841 a_6602_3892.n1 a_6602_3892.n0 172.311
R15842 a_6602_3892.n2 a_6602_3892.n1 24
R15843 a_6602_3892.n1 a_6602_3892.t0 21.212
R15844 a_6615_3907.t0 a_6615_3907.t1 242.857
R15845 a_947_975.n0 a_947_975.t1 358.166
R15846 a_947_975.t4 a_947_975.t5 337.399
R15847 a_947_975.t5 a_947_975.t3 285.986
R15848 a_947_975.n0 a_947_975.t4 282.573
R15849 a_947_975.n1 a_947_975.t0 202.857
R15850 a_947_975.n1 a_947_975.n0 173.817
R15851 a_947_975.n1 a_947_975.t2 20.826
R15852 a_947_975.n2 a_947_975.n1 20.689
R15853 a_3247_4148.n0 a_3247_4148.t0 358.166
R15854 a_3247_4148.t5 a_3247_4148.t3 337.399
R15855 a_3247_4148.t3 a_3247_4148.t4 285.986
R15856 a_3247_4148.n0 a_3247_4148.t5 282.573
R15857 a_3247_4148.n1 a_3247_4148.t2 202.857
R15858 a_3247_4148.n1 a_3247_4148.n0 173.817
R15859 a_3247_4148.n1 a_3247_4148.t1 20.826
R15860 a_3247_4148.n2 a_3247_4148.n1 20.689
R15861 a_3152_4133.n0 a_3152_4133.t1 362.857
R15862 a_3152_4133.t3 a_3152_4133.t4 337.399
R15863 a_3152_4133.t4 a_3152_4133.t5 298.839
R15864 a_3152_4133.n0 a_3152_4133.t3 280.405
R15865 a_3152_4133.n1 a_3152_4133.t2 200
R15866 a_3152_4133.n1 a_3152_4133.n0 172.311
R15867 a_3152_4133.n2 a_3152_4133.n1 24
R15868 a_3152_4133.n1 a_3152_4133.t0 21.212
R15869 a_4397_2180.n0 a_4397_2180.t1 358.166
R15870 a_4397_2180.t5 a_4397_2180.t3 337.399
R15871 a_4397_2180.t3 a_4397_2180.t4 285.986
R15872 a_4397_2180.n0 a_4397_2180.t5 282.573
R15873 a_4397_2180.n1 a_4397_2180.t2 202.857
R15874 a_4397_2180.n1 a_4397_2180.n0 173.817
R15875 a_4397_2180.n1 a_4397_2180.t0 20.826
R15876 a_4397_2180.n2 a_4397_2180.n1 20.689
R15877 a_4302_2165.n0 a_4302_2165.t1 362.857
R15878 a_4302_2165.t5 a_4302_2165.t4 337.399
R15879 a_4302_2165.t4 a_4302_2165.t3 298.839
R15880 a_4302_2165.n0 a_4302_2165.t5 280.405
R15881 a_4302_2165.n1 a_4302_2165.t2 200
R15882 a_4302_2165.n1 a_4302_2165.n0 172.311
R15883 a_4302_2165.n2 a_4302_2165.n1 24
R15884 a_4302_2165.n1 a_4302_2165.t0 21.212
R15885 ADC8_OUT[2].n0 ADC8_OUT[2].t4 1354.27
R15886 ADC8_OUT[2].n0 ADC8_OUT[2].t3 821.954
R15887 ADC8_OUT[2].n3 ADC8_OUT[2].t0 349.397
R15888 ADC8_OUT[2].n2 ADC8_OUT[2].t2 266.575
R15889 ADC8_OUT[2].n1 ADC8_OUT[2].n0 149.035
R15890 ADC8_OUT[2].n1 ADC8_OUT[2].t1 46.723
R15891 ADC8_OUT[2] ADC8_OUT[2].n3 38.029
R15892 ADC8_OUT[2].n3 ADC8_OUT[2].n2 34.635
R15893 ADC8_OUT[2].n2 ADC8_OUT[2].n1 17.317
R15894 a_2108_n953.n25 a_2108_n953.t27 561.971
R15895 a_2108_n953.n0 a_2108_n953.t4 461.908
R15896 a_2108_n953.t12 a_2108_n953.n25 108.635
R15897 a_2108_n953.n0 a_2108_n953.t3 79.512
R15898 a_2108_n953.n24 a_2108_n953.t19 65.401
R15899 a_2108_n953.n23 a_2108_n953.t17 65.401
R15900 a_2108_n953.n22 a_2108_n953.t7 65.401
R15901 a_2108_n953.n21 a_2108_n953.t13 65.401
R15902 a_2108_n953.n20 a_2108_n953.t22 65.401
R15903 a_2108_n953.n19 a_2108_n953.t15 65.401
R15904 a_2108_n953.n18 a_2108_n953.t16 65.401
R15905 a_2108_n953.n17 a_2108_n953.t11 65.401
R15906 a_2108_n953.n16 a_2108_n953.t2 65.401
R15907 a_2108_n953.n15 a_2108_n953.t9 65.401
R15908 a_2108_n953.n14 a_2108_n953.t20 65.401
R15909 a_2108_n953.n13 a_2108_n953.t23 65.401
R15910 a_2108_n953.n12 a_2108_n953.t14 65.401
R15911 a_2108_n953.n11 a_2108_n953.t5 65.401
R15912 a_2108_n953.n10 a_2108_n953.t6 65.401
R15913 a_2108_n953.n9 a_2108_n953.t21 65.401
R15914 a_2108_n953.n8 a_2108_n953.t18 65.401
R15915 a_2108_n953.n7 a_2108_n953.t1 65.401
R15916 a_2108_n953.n6 a_2108_n953.t0 65.401
R15917 a_2108_n953.n5 a_2108_n953.t26 65.401
R15918 a_2108_n953.n4 a_2108_n953.t10 65.401
R15919 a_2108_n953.n3 a_2108_n953.t24 65.401
R15920 a_2108_n953.n2 a_2108_n953.t25 65.401
R15921 a_2108_n953.n1 a_2108_n953.t8 65.401
R15922 a_2108_n953.n1 a_2108_n953.n0 5.64
R15923 a_2108_n953.n25 a_2108_n953.n24 4.438
R15924 a_2108_n953.n23 a_2108_n953.n22 2.524
R15925 a_2108_n953.n3 a_2108_n953.n2 2.498
R15926 a_2108_n953.n17 a_2108_n953.n16 2.364
R15927 a_2108_n953.n9 a_2108_n953.n8 2.355
R15928 a_2108_n953.n2 a_2108_n953.n1 1.998
R15929 a_2108_n953.n4 a_2108_n953.n3 1.998
R15930 a_2108_n953.n5 a_2108_n953.n4 1.998
R15931 a_2108_n953.n6 a_2108_n953.n5 1.998
R15932 a_2108_n953.n7 a_2108_n953.n6 1.998
R15933 a_2108_n953.n8 a_2108_n953.n7 1.998
R15934 a_2108_n953.n10 a_2108_n953.n9 1.998
R15935 a_2108_n953.n11 a_2108_n953.n10 1.998
R15936 a_2108_n953.n12 a_2108_n953.n11 1.998
R15937 a_2108_n953.n13 a_2108_n953.n12 1.998
R15938 a_2108_n953.n14 a_2108_n953.n13 1.998
R15939 a_2108_n953.n15 a_2108_n953.n14 1.998
R15940 a_2108_n953.n16 a_2108_n953.n15 1.998
R15941 a_2108_n953.n18 a_2108_n953.n17 1.998
R15942 a_2108_n953.n19 a_2108_n953.n18 1.998
R15943 a_2108_n953.n20 a_2108_n953.n19 1.998
R15944 a_2108_n953.n21 a_2108_n953.n20 1.998
R15945 a_2108_n953.n22 a_2108_n953.n21 1.998
R15946 a_2108_n953.n24 a_2108_n953.n23 1.998
R15947 a_8422_4445.n0 a_8422_4445.t2 358.166
R15948 a_8422_4445.t5 a_8422_4445.t4 337.399
R15949 a_8422_4445.t4 a_8422_4445.t3 285.986
R15950 a_8422_4445.n0 a_8422_4445.t5 282.573
R15951 a_8422_4445.n1 a_8422_4445.t1 202.857
R15952 a_8422_4445.n1 a_8422_4445.n0 173.817
R15953 a_8422_4445.n1 a_8422_4445.t0 20.826
R15954 a_8422_4445.n2 a_8422_4445.n1 20.689
R15955 a_8792_4445.t0 a_8792_4445.t1 242.857
R15956 RWLB[12].n0 RWLB[12].t7 154.228
R15957 RWLB[12].n14 RWLB[12].t12 149.249
R15958 RWLB[12].n13 RWLB[12].t11 149.249
R15959 RWLB[12].n12 RWLB[12].t3 149.249
R15960 RWLB[12].n11 RWLB[12].t15 149.249
R15961 RWLB[12].n10 RWLB[12].t6 149.249
R15962 RWLB[12].n9 RWLB[12].t5 149.249
R15963 RWLB[12].n8 RWLB[12].t9 149.249
R15964 RWLB[12].n7 RWLB[12].t8 149.249
R15965 RWLB[12].n6 RWLB[12].t1 149.249
R15966 RWLB[12].n5 RWLB[12].t0 149.249
R15967 RWLB[12].n4 RWLB[12].t2 149.249
R15968 RWLB[12].n3 RWLB[12].t13 149.249
R15969 RWLB[12].n2 RWLB[12].t10 149.249
R15970 RWLB[12].n1 RWLB[12].t4 149.249
R15971 RWLB[12].n0 RWLB[12].t14 149.249
R15972 RWLB[12] RWLB[12].n14 47.816
R15973 RWLB[12].n1 RWLB[12].n0 4.979
R15974 RWLB[12].n2 RWLB[12].n1 4.979
R15975 RWLB[12].n3 RWLB[12].n2 4.979
R15976 RWLB[12].n4 RWLB[12].n3 4.979
R15977 RWLB[12].n5 RWLB[12].n4 4.979
R15978 RWLB[12].n6 RWLB[12].n5 4.979
R15979 RWLB[12].n7 RWLB[12].n6 4.979
R15980 RWLB[12].n8 RWLB[12].n7 4.979
R15981 RWLB[12].n9 RWLB[12].n8 4.979
R15982 RWLB[12].n10 RWLB[12].n9 4.979
R15983 RWLB[12].n11 RWLB[12].n10 4.979
R15984 RWLB[12].n12 RWLB[12].n11 4.979
R15985 RWLB[12].n13 RWLB[12].n12 4.979
R15986 RWLB[12].n14 RWLB[12].n13 4.979
R15987 a_5917_693.t0 a_5917_693.t1 242.857
R15988 a_8902_2928.n0 a_8902_2928.t0 362.857
R15989 a_8902_2928.t5 a_8902_2928.t4 337.399
R15990 a_8902_2928.t4 a_8902_2928.t3 298.839
R15991 a_8902_2928.n0 a_8902_2928.t5 280.405
R15992 a_8902_2928.n1 a_8902_2928.t2 200
R15993 a_8902_2928.n1 a_8902_2928.n0 172.311
R15994 a_8902_2928.n2 a_8902_2928.n1 24
R15995 a_8902_2928.n1 a_8902_2928.t1 21.212
R15996 a_8915_2943.t0 a_8915_2943.t1 242.857
R15997 a_3727_1924.n0 a_3727_1924.t1 362.857
R15998 a_3727_1924.t4 a_3727_1924.t5 337.399
R15999 a_3727_1924.t5 a_3727_1924.t3 298.839
R16000 a_3727_1924.n0 a_3727_1924.t4 280.405
R16001 a_3727_1924.n1 a_3727_1924.t0 200
R16002 a_3727_1924.n1 a_3727_1924.n0 172.311
R16003 a_3727_1924.n2 a_3727_1924.n1 24
R16004 a_3727_1924.n1 a_3727_1924.t2 21.212
R16005 a_3740_1939.t0 a_3740_1939.t1 242.857
R16006 a_6027_1924.n0 a_6027_1924.t2 362.857
R16007 a_6027_1924.t3 a_6027_1924.t4 337.399
R16008 a_6027_1924.t4 a_6027_1924.t5 298.839
R16009 a_6027_1924.n0 a_6027_1924.t3 280.405
R16010 a_6027_1924.n1 a_6027_1924.t0 200
R16011 a_6027_1924.n1 a_6027_1924.n0 172.311
R16012 a_6027_1924.n2 a_6027_1924.n1 24
R16013 a_6027_1924.n1 a_6027_1924.t1 21.212
R16014 a_6122_1939.n0 a_6122_1939.t2 358.166
R16015 a_6122_1939.t5 a_6122_1939.t4 337.399
R16016 a_6122_1939.t4 a_6122_1939.t3 285.986
R16017 a_6122_1939.n0 a_6122_1939.t5 282.573
R16018 a_6122_1939.n1 a_6122_1939.t0 202.857
R16019 a_6122_1939.n1 a_6122_1939.n0 173.817
R16020 a_6122_1939.n1 a_6122_1939.t1 20.826
R16021 a_6122_1939.n2 a_6122_1939.n1 20.689
R16022 a_6812_n6503.n0 a_6812_n6503.t1 65.064
R16023 a_6812_n6503.t0 a_6812_n6503.n0 42.011
R16024 a_6812_n6503.n0 a_6812_n6503.t2 2.113
R16025 a_3152_3410.n0 a_3152_3410.t2 362.857
R16026 a_3152_3410.t4 a_3152_3410.t5 337.399
R16027 a_3152_3410.t5 a_3152_3410.t3 298.839
R16028 a_3152_3410.n0 a_3152_3410.t4 280.405
R16029 a_3152_3410.n1 a_3152_3410.t0 200
R16030 a_3152_3410.n1 a_3152_3410.n0 172.311
R16031 a_3152_3410.n2 a_3152_3410.n1 24
R16032 a_3152_3410.n1 a_3152_3410.t1 21.212
R16033 a_3165_3425.t0 a_3165_3425.t1 242.857
R16034 a_4377_n2234.n2 a_4377_n2234.t0 282.97
R16035 a_4377_n2234.n1 a_4377_n2234.t2 240.683
R16036 a_4377_n2234.n0 a_4377_n2234.t3 209.208
R16037 a_4377_n2234.n0 a_4377_n2234.t4 194.167
R16038 a_4377_n2234.t1 a_4377_n2234.n2 183.404
R16039 a_4377_n2234.n1 a_4377_n2234.n0 14.805
R16040 a_4377_n2234.n2 a_4377_n2234.n1 6.415
R16041 a_4618_n2086.t0 a_4618_n2086.t1 34.8
R16042 ADC14_OUT[3].n0 ADC14_OUT[3].t4 1355.37
R16043 ADC14_OUT[3].n0 ADC14_OUT[3].t3 820.859
R16044 ADC14_OUT[3].n3 ADC14_OUT[3].t0 333.655
R16045 ADC14_OUT[3].n2 ADC14_OUT[3].t1 266.644
R16046 ADC14_OUT[3].n1 ADC14_OUT[3].n0 149.035
R16047 ADC14_OUT[3].n3 ADC14_OUT[3].n2 50.447
R16048 ADC14_OUT[3].n1 ADC14_OUT[3].t2 45.968
R16049 ADC14_OUT[3] ADC14_OUT[3].n3 22.133
R16050 ADC14_OUT[3].n2 ADC14_OUT[3].n1 17.317
R16051 a_12963_n8583.n0 a_12963_n8583.t4 1465.51
R16052 a_12963_n8583.n0 a_12963_n8583.t3 712.44
R16053 a_12963_n8583.n1 a_12963_n8583.t0 375.067
R16054 a_12963_n8583.n1 a_12963_n8583.t1 272.668
R16055 a_12963_n8583.n2 a_12963_n8583.n0 143.764
R16056 a_12963_n8583.t2 a_12963_n8583.n2 78.193
R16057 a_12963_n8583.n2 a_12963_n8583.n1 4.517
R16058 a_277_2406.n0 a_277_2406.t1 362.857
R16059 a_277_2406.t5 a_277_2406.t3 337.399
R16060 a_277_2406.t3 a_277_2406.t4 298.839
R16061 a_277_2406.n0 a_277_2406.t5 280.405
R16062 a_277_2406.n1 a_277_2406.t0 200
R16063 a_277_2406.n1 a_277_2406.n0 172.311
R16064 a_277_2406.n2 a_277_2406.n1 24
R16065 a_277_2406.n1 a_277_2406.t2 21.212
R16066 a_372_2421.n0 a_372_2421.t2 358.166
R16067 a_372_2421.t3 a_372_2421.t5 337.399
R16068 a_372_2421.t5 a_372_2421.t4 285.986
R16069 a_372_2421.n0 a_372_2421.t3 282.573
R16070 a_372_2421.n1 a_372_2421.t0 202.857
R16071 a_372_2421.n1 a_372_2421.n0 173.817
R16072 a_372_2421.n1 a_372_2421.t1 20.826
R16073 a_372_2421.n2 a_372_2421.n1 20.689
R16074 a_947_1939.n0 a_947_1939.t0 358.166
R16075 a_947_1939.t4 a_947_1939.t5 337.399
R16076 a_947_1939.t5 a_947_1939.t3 285.986
R16077 a_947_1939.n0 a_947_1939.t4 282.573
R16078 a_947_1939.n1 a_947_1939.t2 202.857
R16079 a_947_1939.n1 a_947_1939.n0 173.817
R16080 a_947_1939.n1 a_947_1939.t1 20.826
R16081 a_947_1939.n2 a_947_1939.n1 20.689
R16082 a_1317_1939.t0 a_1317_1939.t1 242.857
R16083 RWLB[14].n0 RWLB[14].t13 154.228
R16084 RWLB[14].n14 RWLB[14].t2 149.249
R16085 RWLB[14].n13 RWLB[14].t1 149.249
R16086 RWLB[14].n12 RWLB[14].t9 149.249
R16087 RWLB[14].n11 RWLB[14].t5 149.249
R16088 RWLB[14].n10 RWLB[14].t12 149.249
R16089 RWLB[14].n9 RWLB[14].t11 149.249
R16090 RWLB[14].n8 RWLB[14].t15 149.249
R16091 RWLB[14].n7 RWLB[14].t14 149.249
R16092 RWLB[14].n6 RWLB[14].t7 149.249
R16093 RWLB[14].n5 RWLB[14].t6 149.249
R16094 RWLB[14].n4 RWLB[14].t8 149.249
R16095 RWLB[14].n3 RWLB[14].t3 149.249
R16096 RWLB[14].n2 RWLB[14].t0 149.249
R16097 RWLB[14].n1 RWLB[14].t10 149.249
R16098 RWLB[14].n0 RWLB[14].t4 149.249
R16099 RWLB[14] RWLB[14].n14 47.816
R16100 RWLB[14].n1 RWLB[14].n0 4.979
R16101 RWLB[14].n2 RWLB[14].n1 4.979
R16102 RWLB[14].n3 RWLB[14].n2 4.979
R16103 RWLB[14].n4 RWLB[14].n3 4.979
R16104 RWLB[14].n5 RWLB[14].n4 4.979
R16105 RWLB[14].n6 RWLB[14].n5 4.979
R16106 RWLB[14].n7 RWLB[14].n6 4.979
R16107 RWLB[14].n8 RWLB[14].n7 4.979
R16108 RWLB[14].n9 RWLB[14].n8 4.979
R16109 RWLB[14].n10 RWLB[14].n9 4.979
R16110 RWLB[14].n11 RWLB[14].n10 4.979
R16111 RWLB[14].n12 RWLB[14].n11 4.979
R16112 RWLB[14].n13 RWLB[14].n12 4.979
R16113 RWLB[14].n14 RWLB[14].n13 4.979
R16114 a_7642_211.t0 a_7642_211.t1 242.857
R16115 a_6027_678.n0 a_6027_678.t0 362.857
R16116 a_6027_678.t4 a_6027_678.t3 337.399
R16117 a_6027_678.t3 a_6027_678.t5 298.839
R16118 a_6027_678.n0 a_6027_678.t4 280.405
R16119 a_6027_678.n1 a_6027_678.t2 200
R16120 a_6027_678.n1 a_6027_678.n0 172.311
R16121 a_6027_678.n2 a_6027_678.n1 24
R16122 a_6027_678.n1 a_6027_678.t1 21.212
R16123 a_6122_693.n0 a_6122_693.t2 358.166
R16124 a_6122_693.t5 a_6122_693.t4 337.399
R16125 a_6122_693.t4 a_6122_693.t3 285.986
R16126 a_6122_693.n0 a_6122_693.t5 282.573
R16127 a_6122_693.n1 a_6122_693.t0 202.857
R16128 a_6122_693.n1 a_6122_693.n0 173.817
R16129 a_6122_693.n1 a_6122_693.t1 20.826
R16130 a_6122_693.n2 a_6122_693.n1 20.689
R16131 a_13033_n4470.n0 a_13033_n4470.t0 63.08
R16132 a_13033_n4470.n0 a_13033_n4470.t2 41.305
R16133 a_13033_n4470.t1 a_13033_n4470.n0 2.251
R16134 a_13171_n4470.t0 a_13171_n4470.t1 68.741
R16135 a_1522_452.n0 a_1522_452.t1 358.166
R16136 a_1522_452.t3 a_1522_452.t5 337.399
R16137 a_1522_452.t5 a_1522_452.t4 285.986
R16138 a_1522_452.n0 a_1522_452.t3 282.573
R16139 a_1522_452.n1 a_1522_452.t2 202.857
R16140 a_1522_452.n1 a_1522_452.n0 173.817
R16141 a_1522_452.n1 a_1522_452.t0 20.826
R16142 a_1522_452.n2 a_1522_452.n1 20.689
R16143 a_7260_n1770.n0 a_7260_n1770.t2 325.682
R16144 a_7260_n1770.t0 a_7260_n1770.n0 322.293
R16145 a_7260_n1770.n0 a_7260_n1770.t1 73.623
R16146 a_7302_n1770.t0 a_7302_n1770.t1 213.924
R16147 a_7067_n512.t0 a_7067_n512.t1 242.857
R16148 WWLD[5].n0 WWLD[5].t27 262.032
R16149 WWLD[5].n29 WWLD[5].t30 260.715
R16150 WWLD[5].n27 WWLD[5].t0 260.715
R16151 WWLD[5].n25 WWLD[5].t20 260.715
R16152 WWLD[5].n23 WWLD[5].t11 260.715
R16153 WWLD[5].n21 WWLD[5].t22 260.715
R16154 WWLD[5].n19 WWLD[5].t6 260.715
R16155 WWLD[5].n17 WWLD[5].t29 260.715
R16156 WWLD[5].n15 WWLD[5].t16 260.715
R16157 WWLD[5].n13 WWLD[5].t2 260.715
R16158 WWLD[5].n11 WWLD[5].t12 260.715
R16159 WWLD[5].n9 WWLD[5].t31 260.715
R16160 WWLD[5].n7 WWLD[5].t18 260.715
R16161 WWLD[5].n5 WWLD[5].t7 260.715
R16162 WWLD[5].n3 WWLD[5].t23 260.715
R16163 WWLD[5].n1 WWLD[5].t3 260.715
R16164 WWLD[5].n30 WWLD[5].t1 259.254
R16165 WWLD[5].n28 WWLD[5].t10 259.254
R16166 WWLD[5].n26 WWLD[5].t21 259.254
R16167 WWLD[5].n24 WWLD[5].t4 259.254
R16168 WWLD[5].n22 WWLD[5].t26 259.254
R16169 WWLD[5].n20 WWLD[5].t13 259.254
R16170 WWLD[5].n18 WWLD[5].t24 259.254
R16171 WWLD[5].n16 WWLD[5].t8 259.254
R16172 WWLD[5].n14 WWLD[5].t28 259.254
R16173 WWLD[5].n12 WWLD[5].t17 259.254
R16174 WWLD[5].n10 WWLD[5].t5 259.254
R16175 WWLD[5].n8 WWLD[5].t14 259.254
R16176 WWLD[5].n6 WWLD[5].t15 259.254
R16177 WWLD[5].n4 WWLD[5].t19 259.254
R16178 WWLD[5].n2 WWLD[5].t9 259.254
R16179 WWLD[5].n0 WWLD[5].t25 259.254
R16180 WWLD[5] WWLD[5].n30 44.647
R16181 WWLD[5].n1 WWLD[5].n0 3.576
R16182 WWLD[5].n3 WWLD[5].n2 3.576
R16183 WWLD[5].n5 WWLD[5].n4 3.576
R16184 WWLD[5].n7 WWLD[5].n6 3.576
R16185 WWLD[5].n9 WWLD[5].n8 3.576
R16186 WWLD[5].n11 WWLD[5].n10 3.576
R16187 WWLD[5].n13 WWLD[5].n12 3.576
R16188 WWLD[5].n15 WWLD[5].n14 3.576
R16189 WWLD[5].n17 WWLD[5].n16 3.576
R16190 WWLD[5].n19 WWLD[5].n18 3.576
R16191 WWLD[5].n21 WWLD[5].n20 3.576
R16192 WWLD[5].n23 WWLD[5].n22 3.576
R16193 WWLD[5].n25 WWLD[5].n24 3.576
R16194 WWLD[5].n27 WWLD[5].n26 3.576
R16195 WWLD[5].n29 WWLD[5].n28 3.576
R16196 WWLD[5].n2 WWLD[5].n1 1.317
R16197 WWLD[5].n4 WWLD[5].n3 1.317
R16198 WWLD[5].n6 WWLD[5].n5 1.317
R16199 WWLD[5].n8 WWLD[5].n7 1.317
R16200 WWLD[5].n10 WWLD[5].n9 1.317
R16201 WWLD[5].n12 WWLD[5].n11 1.317
R16202 WWLD[5].n14 WWLD[5].n13 1.317
R16203 WWLD[5].n16 WWLD[5].n15 1.317
R16204 WWLD[5].n18 WWLD[5].n17 1.317
R16205 WWLD[5].n20 WWLD[5].n19 1.317
R16206 WWLD[5].n22 WWLD[5].n21 1.317
R16207 WWLD[5].n24 WWLD[5].n23 1.317
R16208 WWLD[5].n26 WWLD[5].n25 1.317
R16209 WWLD[5].n28 WWLD[5].n27 1.317
R16210 WWLD[5].n30 WWLD[5].n29 1.317
R16211 a_852_n527.n0 a_852_n527.t1 362.857
R16212 a_852_n527.t3 a_852_n527.t4 337.399
R16213 a_852_n527.t4 a_852_n527.t5 298.839
R16214 a_852_n527.n0 a_852_n527.t3 280.405
R16215 a_852_n527.n1 a_852_n527.t0 200
R16216 a_852_n527.n1 a_852_n527.n0 172.311
R16217 a_852_n527.n2 a_852_n527.n1 24
R16218 a_852_n527.n1 a_852_n527.t2 21.212
R16219 ADC1_OUT[2].n0 ADC1_OUT[2].t4 1354.27
R16220 ADC1_OUT[2].n0 ADC1_OUT[2].t3 821.954
R16221 ADC1_OUT[2].n3 ADC1_OUT[2].t0 347.891
R16222 ADC1_OUT[2].n2 ADC1_OUT[2].t1 266.575
R16223 ADC1_OUT[2].n1 ADC1_OUT[2].n0 149.035
R16224 ADC1_OUT[2].n1 ADC1_OUT[2].t2 46.723
R16225 ADC1_OUT[2] ADC1_OUT[2].n3 38.02
R16226 ADC1_OUT[2].n3 ADC1_OUT[2].n2 36.141
R16227 ADC1_OUT[2].n2 ADC1_OUT[2].n1 17.317
R16228 a_8935_n1371.n1 a_8935_n1371.t4 550.94
R16229 a_8935_n1371.n1 a_8935_n1371.t3 500.621
R16230 a_8935_n1371.t2 a_8935_n1371.n2 192.787
R16231 a_8935_n1371.n0 a_8935_n1371.t0 163.997
R16232 a_8935_n1371.n2 a_8935_n1371.n1 149.035
R16233 a_8935_n1371.n0 a_8935_n1371.t1 54.068
R16234 a_8935_n1371.n2 a_8935_n1371.n0 17.317
R16235 a_7847_4686.n0 a_7847_4686.t1 358.166
R16236 a_7847_4686.t5 a_7847_4686.t3 337.399
R16237 a_7847_4686.t3 a_7847_4686.t4 285.986
R16238 a_7847_4686.n0 a_7847_4686.t5 282.573
R16239 a_7847_4686.n1 a_7847_4686.t2 202.857
R16240 a_7847_4686.n1 a_7847_4686.n0 173.817
R16241 a_7847_4686.n1 a_7847_4686.t0 20.826
R16242 a_7847_4686.n2 a_7847_4686.n1 20.689
R16243 a_4302_3892.n0 a_4302_3892.t1 362.857
R16244 a_4302_3892.t4 a_4302_3892.t3 337.399
R16245 a_4302_3892.t3 a_4302_3892.t5 298.839
R16246 a_4302_3892.n0 a_4302_3892.t4 280.405
R16247 a_4302_3892.n1 a_4302_3892.t0 200
R16248 a_4302_3892.n1 a_4302_3892.n0 172.311
R16249 a_4302_3892.n2 a_4302_3892.n1 24
R16250 a_4302_3892.n1 a_4302_3892.t2 21.212
R16251 a_4397_3907.n0 a_4397_3907.t1 358.166
R16252 a_4397_3907.t4 a_4397_3907.t5 337.399
R16253 a_4397_3907.t5 a_4397_3907.t3 285.986
R16254 a_4397_3907.n0 a_4397_3907.t4 282.573
R16255 a_4397_3907.n1 a_4397_3907.t2 202.857
R16256 a_4397_3907.n1 a_4397_3907.n0 173.817
R16257 a_4397_3907.n1 a_4397_3907.t0 20.826
R16258 a_4397_3907.n2 a_4397_3907.n1 20.689
R16259 a_1427_1442.n0 a_1427_1442.t1 362.857
R16260 a_1427_1442.t5 a_1427_1442.t3 337.399
R16261 a_1427_1442.t3 a_1427_1442.t4 298.839
R16262 a_1427_1442.n0 a_1427_1442.t5 280.405
R16263 a_1427_1442.n1 a_1427_1442.t2 200
R16264 a_1427_1442.n1 a_1427_1442.n0 172.311
R16265 a_1427_1442.n2 a_1427_1442.n1 24
R16266 a_1427_1442.n1 a_1427_1442.t0 21.212
R16267 a_1522_1457.n0 a_1522_1457.t1 358.166
R16268 a_1522_1457.t4 a_1522_1457.t3 337.399
R16269 a_1522_1457.t3 a_1522_1457.t5 285.986
R16270 a_1522_1457.n0 a_1522_1457.t4 282.573
R16271 a_1522_1457.n1 a_1522_1457.t2 202.857
R16272 a_1522_1457.n1 a_1522_1457.n0 173.817
R16273 a_1522_1457.n1 a_1522_1457.t0 20.826
R16274 a_1522_1457.n2 a_1522_1457.n1 20.689
R16275 a_7190_4148.t0 a_7190_4148.t1 242.857
R16276 a_8327_3651.n0 a_8327_3651.t1 362.857
R16277 a_8327_3651.t3 a_8327_3651.t4 337.399
R16278 a_8327_3651.t4 a_8327_3651.t5 298.839
R16279 a_8327_3651.n0 a_8327_3651.t3 280.405
R16280 a_8327_3651.n1 a_8327_3651.t2 200
R16281 a_8327_3651.n1 a_8327_3651.n0 172.311
R16282 a_8327_3651.n2 a_8327_3651.n1 24
R16283 a_8327_3651.n1 a_8327_3651.t0 21.212
R16284 a_8422_3666.n0 a_8422_3666.t1 358.166
R16285 a_8422_3666.t5 a_8422_3666.t4 337.399
R16286 a_8422_3666.t4 a_8422_3666.t3 285.986
R16287 a_8422_3666.n0 a_8422_3666.t5 282.573
R16288 a_8422_3666.n1 a_8422_3666.t2 202.857
R16289 a_8422_3666.n1 a_8422_3666.n0 173.817
R16290 a_8422_3666.n1 a_8422_3666.t0 20.826
R16291 a_8422_3666.n2 a_8422_3666.n1 20.689
R16292 a_n2415_n5850.n0 a_n2415_n5850.t3 1465.51
R16293 a_n2415_n5850.n0 a_n2415_n5850.t4 712.44
R16294 a_n2415_n5850.n1 a_n2415_n5850.t0 375.067
R16295 a_n2415_n5850.n1 a_n2415_n5850.t1 272.668
R16296 a_n2415_n5850.n2 a_n2415_n5850.n0 143.764
R16297 a_n2415_n5850.t2 a_n2415_n5850.n2 78.193
R16298 a_n2415_n5850.n2 a_n2415_n5850.n1 4.517
R16299 a_6602_2928.n0 a_6602_2928.t1 362.857
R16300 a_6602_2928.t4 a_6602_2928.t3 337.399
R16301 a_6602_2928.t3 a_6602_2928.t5 298.839
R16302 a_6602_2928.n0 a_6602_2928.t4 280.405
R16303 a_6602_2928.n1 a_6602_2928.t2 200
R16304 a_6602_2928.n1 a_6602_2928.n0 172.311
R16305 a_6602_2928.n2 a_6602_2928.n1 24
R16306 a_6602_2928.n1 a_6602_2928.t0 21.212
R16307 a_6697_2943.n0 a_6697_2943.t2 358.166
R16308 a_6697_2943.t4 a_6697_2943.t5 337.399
R16309 a_6697_2943.t5 a_6697_2943.t3 285.986
R16310 a_6697_2943.n0 a_6697_2943.t4 282.573
R16311 a_6697_2943.n1 a_6697_2943.t0 202.857
R16312 a_6697_2943.n1 a_6697_2943.n0 173.817
R16313 a_6697_2943.n1 a_6697_2943.t1 20.826
R16314 a_6697_2943.n2 a_6697_2943.n1 20.689
R16315 RWLB[8].n0 RWLB[8].t13 154.228
R16316 RWLB[8].n14 RWLB[8].t14 149.249
R16317 RWLB[8].n13 RWLB[8].t0 149.249
R16318 RWLB[8].n12 RWLB[8].t11 149.249
R16319 RWLB[8].n11 RWLB[8].t5 149.249
R16320 RWLB[8].n10 RWLB[8].t15 149.249
R16321 RWLB[8].n9 RWLB[8].t2 149.249
R16322 RWLB[8].n8 RWLB[8].t3 149.249
R16323 RWLB[8].n7 RWLB[8].t8 149.249
R16324 RWLB[8].n6 RWLB[8].t1 149.249
R16325 RWLB[8].n5 RWLB[8].t6 149.249
R16326 RWLB[8].n4 RWLB[8].t7 149.249
R16327 RWLB[8].n3 RWLB[8].t12 149.249
R16328 RWLB[8].n2 RWLB[8].t4 149.249
R16329 RWLB[8].n1 RWLB[8].t10 149.249
R16330 RWLB[8].n0 RWLB[8].t9 149.249
R16331 RWLB[8] RWLB[8].n14 47.816
R16332 RWLB[8].n1 RWLB[8].n0 4.979
R16333 RWLB[8].n2 RWLB[8].n1 4.979
R16334 RWLB[8].n3 RWLB[8].n2 4.979
R16335 RWLB[8].n4 RWLB[8].n3 4.979
R16336 RWLB[8].n5 RWLB[8].n4 4.979
R16337 RWLB[8].n6 RWLB[8].n5 4.979
R16338 RWLB[8].n7 RWLB[8].n6 4.979
R16339 RWLB[8].n8 RWLB[8].n7 4.979
R16340 RWLB[8].n9 RWLB[8].n8 4.979
R16341 RWLB[8].n10 RWLB[8].n9 4.979
R16342 RWLB[8].n11 RWLB[8].n10 4.979
R16343 RWLB[8].n12 RWLB[8].n11 4.979
R16344 RWLB[8].n13 RWLB[8].n12 4.979
R16345 RWLB[8].n14 RWLB[8].n13 4.979
R16346 a_1317_1698.t0 a_1317_1698.t1 242.857
R16347 a_6492_693.t0 a_6492_693.t1 242.857
R16348 ADC6_OUT[1].n0 ADC6_OUT[1].t3 1355.37
R16349 ADC6_OUT[1].n0 ADC6_OUT[1].t4 820.859
R16350 ADC6_OUT[1].n3 ADC6_OUT[1].t0 338.173
R16351 ADC6_OUT[1].n2 ADC6_OUT[1].t1 266.644
R16352 ADC6_OUT[1].n1 ADC6_OUT[1].n0 149.035
R16353 ADC6_OUT[1].n1 ADC6_OUT[1].t2 45.968
R16354 ADC6_OUT[1].n3 ADC6_OUT[1].n2 45.929
R16355 ADC6_OUT[1] ADC6_OUT[1].n3 45.856
R16356 ADC6_OUT[1].n2 ADC6_OUT[1].n1 17.317
R16357 a_3563_n5338.n0 a_3563_n5338.t0 63.08
R16358 a_3563_n5338.n0 a_3563_n5338.t2 41.307
R16359 a_3563_n5338.t1 a_3563_n5338.n0 2.251
R16360 a_3493_n5850.n0 a_3493_n5850.t4 1465.51
R16361 a_3493_n5850.n0 a_3493_n5850.t3 712.44
R16362 a_3493_n5850.n1 a_3493_n5850.t0 375.067
R16363 a_3493_n5850.n1 a_3493_n5850.t2 272.668
R16364 a_3493_n5850.n2 a_3493_n5850.n0 143.764
R16365 a_3493_n5850.t1 a_3493_n5850.n2 78.193
R16366 a_3493_n5850.n2 a_3493_n5850.n1 4.517
R16367 a_4972_n30.n0 a_4972_n30.t1 358.166
R16368 a_4972_n30.t5 a_4972_n30.t3 337.399
R16369 a_4972_n30.t3 a_4972_n30.t4 285.986
R16370 a_4972_n30.n0 a_4972_n30.t5 282.573
R16371 a_4972_n30.n1 a_4972_n30.t2 202.857
R16372 a_4972_n30.n1 a_4972_n30.n0 173.817
R16373 a_4972_n30.n1 a_4972_n30.t0 20.826
R16374 a_4972_n30.n2 a_4972_n30.n1 20.689
R16375 a_4877_n45.n0 a_4877_n45.t1 362.857
R16376 a_4877_n45.t4 a_4877_n45.t3 337.399
R16377 a_4877_n45.t3 a_4877_n45.t5 298.839
R16378 a_4877_n45.n0 a_4877_n45.t4 280.405
R16379 a_4877_n45.n1 a_4877_n45.t2 200
R16380 a_4877_n45.n1 a_4877_n45.n0 172.311
R16381 a_4877_n45.n2 a_4877_n45.n1 24
R16382 a_4877_n45.n1 a_4877_n45.t0 21.212
R16383 a_2015_211.t0 a_2015_211.t1 242.857
R16384 PRE_A.n14 PRE_A.t14 334.341
R16385 PRE_A.n7 PRE_A.t6 330.621
R16386 PRE_A.n8 PRE_A.t1 330.576
R16387 PRE_A.n10 PRE_A.t7 330.576
R16388 PRE_A.n1 PRE_A.t13 329.868
R16389 PRE_A.n0 PRE_A.t3 329.823
R16390 PRE_A.n13 PRE_A.t11 329.115
R16391 PRE_A.n2 PRE_A.t10 329.07
R16392 PRE_A.n11 PRE_A.t12 328.362
R16393 PRE_A.n3 PRE_A.t2 327.609
R16394 PRE_A.n5 PRE_A.t0 327.609
R16395 PRE_A.n9 PRE_A.t4 327.609
R16396 PRE_A.n6 PRE_A.t15 327.564
R16397 PRE_A.n4 PRE_A.t8 326.058
R16398 PRE_A.n12 PRE_A.t5 326.058
R16399 PRE_A.n0 PRE_A.t9 315.213
R16400 PRE_A PRE_A.n14 7.853
R16401 PRE_A.n6 PRE_A.n5 1.072
R16402 PRE_A.n14 PRE_A.n13 1.071
R16403 PRE_A.n12 PRE_A.n11 1.07
R16404 PRE_A.n2 PRE_A.n1 1.07
R16405 PRE_A.n10 PRE_A.n9 1.07
R16406 PRE_A.n4 PRE_A.n3 1.068
R16407 PRE_A.n8 PRE_A.n7 1.068
R16408 PRE_A.n11 PRE_A.n10 0.705
R16409 PRE_A.n1 PRE_A.n0 0.703
R16410 PRE_A.n3 PRE_A.n2 0.703
R16411 PRE_A.n7 PRE_A.n6 0.703
R16412 PRE_A.n9 PRE_A.n8 0.703
R16413 PRE_A.n5 PRE_A.n4 0.7
R16414 PRE_A.n13 PRE_A.n12 0.697
R16415 a_5543_n2422.n3 a_5543_n2422.t1 475.39
R16416 a_5543_n2422.n3 a_5543_n2422.n2 422.502
R16417 a_5543_n2422.t4 a_5543_n2422.t6 228.696
R16418 a_5543_n2422.n2 a_5543_n2422.t3 185.704
R16419 a_5543_n2422.n0 a_5543_n2422.t4 126.761
R16420 a_5543_n2422.n1 a_5543_n2422.t5 126.284
R16421 a_5543_n2422.n1 a_5543_n2422.t2 126.284
R16422 a_5543_n2422.t0 a_5543_n2422.n3 124.375
R16423 a_5543_n2422.t2 a_5543_n2422.n0 115.122
R16424 a_5543_n2422.n0 a_5543_n2422.t7 111.229
R16425 a_5543_n2422.n2 a_5543_n2422.n1 8.764
R16426 a_1427_960.n0 a_1427_960.t2 362.857
R16427 a_1427_960.t3 a_1427_960.t5 337.399
R16428 a_1427_960.t5 a_1427_960.t4 298.839
R16429 a_1427_960.n0 a_1427_960.t3 280.405
R16430 a_1427_960.n1 a_1427_960.t0 200
R16431 a_1427_960.n1 a_1427_960.n0 172.311
R16432 a_1427_960.n2 a_1427_960.n1 24
R16433 a_1427_960.n1 a_1427_960.t1 21.212
R16434 a_1522_975.n0 a_1522_975.t2 358.166
R16435 a_1522_975.t5 a_1522_975.t4 337.399
R16436 a_1522_975.t4 a_1522_975.t3 285.986
R16437 a_1522_975.n0 a_1522_975.t5 282.573
R16438 a_1522_975.n1 a_1522_975.t0 202.857
R16439 a_1522_975.n1 a_1522_975.n0 173.817
R16440 a_1522_975.n1 a_1522_975.t1 20.826
R16441 a_1522_975.n2 a_1522_975.n1 20.689
R16442 a_9143_n6849.t1 a_9143_n6849.t0 42.707
R16443 a_9178_n6503.n0 a_9178_n6503.t0 65.064
R16444 a_9178_n6503.t1 a_9178_n6503.n0 42.011
R16445 a_9178_n6503.n0 a_9178_n6503.t2 2.113
R16446 a_6122_3184.n0 a_6122_3184.t2 358.166
R16447 a_6122_3184.t5 a_6122_3184.t4 337.399
R16448 a_6122_3184.t4 a_6122_3184.t3 285.986
R16449 a_6122_3184.n0 a_6122_3184.t5 282.573
R16450 a_6122_3184.n1 a_6122_3184.t1 202.857
R16451 a_6122_3184.n1 a_6122_3184.n0 173.817
R16452 a_6122_3184.n1 a_6122_3184.t0 20.826
R16453 a_6122_3184.n2 a_6122_3184.n1 20.689
R16454 a_6492_3184.t0 a_6492_3184.t1 242.857
R16455 WWL[5].n0 WWL[5].t15 262.032
R16456 WWL[5].n29 WWL[5].t18 260.715
R16457 WWL[5].n27 WWL[5].t21 260.715
R16458 WWL[5].n25 WWL[5].t3 260.715
R16459 WWL[5].n23 WWL[5].t29 260.715
R16460 WWL[5].n21 WWL[5].t9 260.715
R16461 WWL[5].n19 WWL[5].t26 260.715
R16462 WWL[5].n17 WWL[5].t17 260.715
R16463 WWL[5].n15 WWL[5].t0 260.715
R16464 WWL[5].n13 WWL[5].t22 260.715
R16465 WWL[5].n11 WWL[5].t30 260.715
R16466 WWL[5].n9 WWL[5].t19 260.715
R16467 WWL[5].n7 WWL[5].t1 260.715
R16468 WWL[5].n5 WWL[5].t27 260.715
R16469 WWL[5].n3 WWL[5].t10 260.715
R16470 WWL[5].n1 WWL[5].t23 260.715
R16471 WWL[5].n30 WWL[5].t2 259.254
R16472 WWL[5].n28 WWL[5].t8 259.254
R16473 WWL[5].n26 WWL[5].t20 259.254
R16474 WWL[5].n24 WWL[5].t4 259.254
R16475 WWL[5].n22 WWL[5].t28 259.254
R16476 WWL[5].n20 WWL[5].t11 259.254
R16477 WWL[5].n18 WWL[5].t24 259.254
R16478 WWL[5].n16 WWL[5].t6 259.254
R16479 WWL[5].n14 WWL[5].t31 259.254
R16480 WWL[5].n12 WWL[5].t14 259.254
R16481 WWL[5].n10 WWL[5].t5 259.254
R16482 WWL[5].n8 WWL[5].t12 259.254
R16483 WWL[5].n6 WWL[5].t13 259.254
R16484 WWL[5].n4 WWL[5].t16 259.254
R16485 WWL[5].n2 WWL[5].t7 259.254
R16486 WWL[5].n0 WWL[5].t25 259.254
R16487 WWL[5] WWL[5].n30 44.647
R16488 WWL[5].n1 WWL[5].n0 3.576
R16489 WWL[5].n3 WWL[5].n2 3.576
R16490 WWL[5].n5 WWL[5].n4 3.576
R16491 WWL[5].n7 WWL[5].n6 3.576
R16492 WWL[5].n9 WWL[5].n8 3.576
R16493 WWL[5].n11 WWL[5].n10 3.576
R16494 WWL[5].n13 WWL[5].n12 3.576
R16495 WWL[5].n15 WWL[5].n14 3.576
R16496 WWL[5].n17 WWL[5].n16 3.576
R16497 WWL[5].n19 WWL[5].n18 3.576
R16498 WWL[5].n21 WWL[5].n20 3.576
R16499 WWL[5].n23 WWL[5].n22 3.576
R16500 WWL[5].n25 WWL[5].n24 3.576
R16501 WWL[5].n27 WWL[5].n26 3.576
R16502 WWL[5].n29 WWL[5].n28 3.576
R16503 WWL[5].n2 WWL[5].n1 1.317
R16504 WWL[5].n4 WWL[5].n3 1.317
R16505 WWL[5].n6 WWL[5].n5 1.317
R16506 WWL[5].n8 WWL[5].n7 1.317
R16507 WWL[5].n10 WWL[5].n9 1.317
R16508 WWL[5].n12 WWL[5].n11 1.317
R16509 WWL[5].n14 WWL[5].n13 1.317
R16510 WWL[5].n16 WWL[5].n15 1.317
R16511 WWL[5].n18 WWL[5].n17 1.317
R16512 WWL[5].n20 WWL[5].n19 1.317
R16513 WWL[5].n22 WWL[5].n21 1.317
R16514 WWL[5].n24 WWL[5].n23 1.317
R16515 WWL[5].n26 WWL[5].n25 1.317
R16516 WWL[5].n28 WWL[5].n27 1.317
R16517 WWL[5].n30 WWL[5].n29 1.317
R16518 a_4302_2406.n0 a_4302_2406.t2 362.857
R16519 a_4302_2406.t3 a_4302_2406.t5 337.399
R16520 a_4302_2406.t5 a_4302_2406.t4 298.839
R16521 a_4302_2406.n0 a_4302_2406.t3 280.405
R16522 a_4302_2406.n1 a_4302_2406.t1 200
R16523 a_4302_2406.n1 a_4302_2406.n0 172.311
R16524 a_4302_2406.n2 a_4302_2406.n1 24
R16525 a_4302_2406.n1 a_4302_2406.t0 21.212
R16526 a_7177_437.n0 a_7177_437.t2 362.857
R16527 a_7177_437.t3 a_7177_437.t5 337.399
R16528 a_7177_437.t5 a_7177_437.t4 298.839
R16529 a_7177_437.n0 a_7177_437.t3 280.405
R16530 a_7177_437.n1 a_7177_437.t1 200
R16531 a_7177_437.n1 a_7177_437.n0 172.311
R16532 a_7177_437.n2 a_7177_437.n1 24
R16533 a_7177_437.n1 a_7177_437.t0 21.212
R16534 a_7272_452.n0 a_7272_452.t2 358.166
R16535 a_7272_452.t4 a_7272_452.t3 337.399
R16536 a_7272_452.t3 a_7272_452.t5 285.986
R16537 a_7272_452.n0 a_7272_452.t4 282.573
R16538 a_7272_452.n1 a_7272_452.t0 202.857
R16539 a_7272_452.n1 a_7272_452.n0 173.817
R16540 a_7272_452.n1 a_7272_452.t1 20.826
R16541 a_7272_452.n2 a_7272_452.n1 20.689
R16542 a_852_196.n0 a_852_196.t2 362.857
R16543 a_852_196.t4 a_852_196.t3 337.399
R16544 a_852_196.t3 a_852_196.t5 298.839
R16545 a_852_196.n0 a_852_196.t4 280.405
R16546 a_852_196.n1 a_852_196.t0 200
R16547 a_852_196.n1 a_852_196.n0 172.311
R16548 a_852_196.n2 a_852_196.n1 24
R16549 a_852_196.n1 a_852_196.t1 21.212
R16550 a_5558_n953.n25 a_5558_n953.t27 561.971
R16551 a_5558_n953.n0 a_5558_n953.t3 461.908
R16552 a_5558_n953.t12 a_5558_n953.n25 108.635
R16553 a_5558_n953.n0 a_5558_n953.t4 79.512
R16554 a_5558_n953.n24 a_5558_n953.t19 65.401
R16555 a_5558_n953.n23 a_5558_n953.t17 65.401
R16556 a_5558_n953.n22 a_5558_n953.t11 65.401
R16557 a_5558_n953.n21 a_5558_n953.t13 65.401
R16558 a_5558_n953.n20 a_5558_n953.t22 65.401
R16559 a_5558_n953.n19 a_5558_n953.t15 65.401
R16560 a_5558_n953.n18 a_5558_n953.t16 65.401
R16561 a_5558_n953.n17 a_5558_n953.t9 65.401
R16562 a_5558_n953.n16 a_5558_n953.t2 65.401
R16563 a_5558_n953.n15 a_5558_n953.t7 65.401
R16564 a_5558_n953.n14 a_5558_n953.t20 65.401
R16565 a_5558_n953.n13 a_5558_n953.t5 65.401
R16566 a_5558_n953.n12 a_5558_n953.t14 65.401
R16567 a_5558_n953.n11 a_5558_n953.t25 65.401
R16568 a_5558_n953.n10 a_5558_n953.t10 65.401
R16569 a_5558_n953.n9 a_5558_n953.t21 65.401
R16570 a_5558_n953.n8 a_5558_n953.t18 65.401
R16571 a_5558_n953.n7 a_5558_n953.t1 65.401
R16572 a_5558_n953.n6 a_5558_n953.t0 65.401
R16573 a_5558_n953.n5 a_5558_n953.t26 65.401
R16574 a_5558_n953.n4 a_5558_n953.t8 65.401
R16575 a_5558_n953.n3 a_5558_n953.t23 65.401
R16576 a_5558_n953.n2 a_5558_n953.t24 65.401
R16577 a_5558_n953.n1 a_5558_n953.t6 65.401
R16578 a_5558_n953.n1 a_5558_n953.n0 5.64
R16579 a_5558_n953.n25 a_5558_n953.n24 4.438
R16580 a_5558_n953.n23 a_5558_n953.n22 2.524
R16581 a_5558_n953.n3 a_5558_n953.n2 2.498
R16582 a_5558_n953.n17 a_5558_n953.n16 2.364
R16583 a_5558_n953.n9 a_5558_n953.n8 2.355
R16584 a_5558_n953.n2 a_5558_n953.n1 1.998
R16585 a_5558_n953.n4 a_5558_n953.n3 1.998
R16586 a_5558_n953.n5 a_5558_n953.n4 1.998
R16587 a_5558_n953.n6 a_5558_n953.n5 1.998
R16588 a_5558_n953.n7 a_5558_n953.n6 1.998
R16589 a_5558_n953.n8 a_5558_n953.n7 1.998
R16590 a_5558_n953.n10 a_5558_n953.n9 1.998
R16591 a_5558_n953.n11 a_5558_n953.n10 1.998
R16592 a_5558_n953.n12 a_5558_n953.n11 1.998
R16593 a_5558_n953.n13 a_5558_n953.n12 1.998
R16594 a_5558_n953.n14 a_5558_n953.n13 1.998
R16595 a_5558_n953.n15 a_5558_n953.n14 1.998
R16596 a_5558_n953.n16 a_5558_n953.n15 1.998
R16597 a_5558_n953.n18 a_5558_n953.n17 1.998
R16598 a_5558_n953.n19 a_5558_n953.n18 1.998
R16599 a_5558_n953.n20 a_5558_n953.n19 1.998
R16600 a_5558_n953.n21 a_5558_n953.n20 1.998
R16601 a_5558_n953.n22 a_5558_n953.n21 1.998
R16602 a_5558_n953.n24 a_5558_n953.n23 1.998
R16603 a_7177_3892.n0 a_7177_3892.t2 362.857
R16604 a_7177_3892.t4 a_7177_3892.t5 337.399
R16605 a_7177_3892.t5 a_7177_3892.t3 298.839
R16606 a_7177_3892.n0 a_7177_3892.t4 280.405
R16607 a_7177_3892.n1 a_7177_3892.t0 200
R16608 a_7177_3892.n1 a_7177_3892.n0 172.311
R16609 a_7177_3892.n2 a_7177_3892.n1 24
R16610 a_7177_3892.n1 a_7177_3892.t1 21.212
R16611 a_7190_3907.t0 a_7190_3907.t1 242.857
R16612 a_6615_3425.t0 a_6615_3425.t1 242.857
R16613 a_8340_2421.t0 a_8340_2421.t1 242.857
R16614 a_7752_1442.n0 a_7752_1442.t2 362.857
R16615 a_7752_1442.t4 a_7752_1442.t5 337.399
R16616 a_7752_1442.t5 a_7752_1442.t3 298.839
R16617 a_7752_1442.n0 a_7752_1442.t4 280.405
R16618 a_7752_1442.n1 a_7752_1442.t0 200
R16619 a_7752_1442.n1 a_7752_1442.n0 172.311
R16620 a_7752_1442.n2 a_7752_1442.n1 24
R16621 a_7752_1442.n1 a_7752_1442.t1 21.212
R16622 a_7765_1457.t0 a_7765_1457.t1 242.857
R16623 a_4302_n286.n0 a_4302_n286.t2 362.857
R16624 a_4302_n286.t3 a_4302_n286.t5 337.399
R16625 a_4302_n286.t5 a_4302_n286.t4 298.839
R16626 a_4302_n286.n0 a_4302_n286.t3 280.405
R16627 a_4302_n286.n1 a_4302_n286.t1 200
R16628 a_4302_n286.n1 a_4302_n286.n0 172.311
R16629 a_4302_n286.n2 a_4302_n286.n1 24
R16630 a_4302_n286.n1 a_4302_n286.t0 21.212
R16631 a_4942_n8026.t1 a_4942_n8026.t0 336.814
R16632 a_4883_n8071.t0 a_4883_n8071.t1 68.74
R16633 a_3822_4148.n0 a_3822_4148.t0 358.166
R16634 a_3822_4148.t4 a_3822_4148.t3 337.399
R16635 a_3822_4148.t3 a_3822_4148.t5 285.986
R16636 a_3822_4148.n0 a_3822_4148.t4 282.573
R16637 a_3822_4148.n1 a_3822_4148.t2 202.857
R16638 a_3822_4148.n1 a_3822_4148.n0 173.817
R16639 a_3822_4148.n1 a_3822_4148.t1 20.826
R16640 a_3822_4148.n2 a_3822_4148.n1 20.689
R16641 a_3727_4133.n0 a_3727_4133.t1 362.857
R16642 a_3727_4133.t3 a_3727_4133.t4 337.399
R16643 a_3727_4133.t4 a_3727_4133.t5 298.839
R16644 a_3727_4133.n0 a_3727_4133.t3 280.405
R16645 a_3727_4133.n1 a_3727_4133.t2 200
R16646 a_3727_4133.n1 a_3727_4133.n0 172.311
R16647 a_3727_4133.n2 a_3727_4133.n1 24
R16648 a_3727_4133.n1 a_3727_4133.t0 21.212
R16649 a_3740_211.t0 a_3740_211.t1 242.857
R16650 a_n52_n7216.n0 a_n52_n7216.t3 1464.36
R16651 a_n52_n7216.n0 a_n52_n7216.t4 713.588
R16652 a_n52_n7216.n1 a_n52_n7216.t0 374.998
R16653 a_n52_n7216.n1 a_n52_n7216.t1 273.351
R16654 a_n52_n7216.n2 a_n52_n7216.n0 143.764
R16655 a_n52_n7216.t2 a_n52_n7216.n2 78.209
R16656 a_n52_n7216.n2 a_n52_n7216.n1 4.517
R16657 ADC3_OUT[2].n0 ADC3_OUT[2].t4 1354.27
R16658 ADC3_OUT[2].n0 ADC3_OUT[2].t3 821.954
R16659 ADC3_OUT[2].n3 ADC3_OUT[2].t0 342.621
R16660 ADC3_OUT[2].n2 ADC3_OUT[2].t2 266.575
R16661 ADC3_OUT[2].n1 ADC3_OUT[2].n0 149.035
R16662 ADC3_OUT[2].n1 ADC3_OUT[2].t1 46.723
R16663 ADC3_OUT[2].n3 ADC3_OUT[2].n2 41.411
R16664 ADC3_OUT[2] ADC3_OUT[2].n3 37.764
R16665 ADC3_OUT[2].n2 ADC3_OUT[2].n1 17.317
R16666 a_n279_n6503.n0 a_n279_n6503.t0 65.064
R16667 a_n279_n6503.n0 a_n279_n6503.t2 42.011
R16668 a_n279_n6503.t1 a_n279_n6503.n0 2.113
R16669 a_865_2421.t0 a_865_2421.t1 242.857
R16670 a_4397_2421.n0 a_4397_2421.t2 358.166
R16671 a_4397_2421.t4 a_4397_2421.t5 337.399
R16672 a_4397_2421.t5 a_4397_2421.t3 285.986
R16673 a_4397_2421.n0 a_4397_2421.t4 282.573
R16674 a_4397_2421.n1 a_4397_2421.t0 202.857
R16675 a_4397_2421.n1 a_4397_2421.n0 173.817
R16676 a_4397_2421.n1 a_4397_2421.t1 20.826
R16677 a_4397_2421.n2 a_4397_2421.n1 20.689
R16678 a_4767_2421.t0 a_4767_2421.t1 242.857
R16679 a_2672_211.n0 a_2672_211.t2 358.166
R16680 a_2672_211.t4 a_2672_211.t3 337.399
R16681 a_2672_211.t3 a_2672_211.t5 285.986
R16682 a_2672_211.n0 a_2672_211.t4 282.573
R16683 a_2672_211.n1 a_2672_211.t1 202.857
R16684 a_2672_211.n1 a_2672_211.n0 173.817
R16685 a_2672_211.n1 a_2672_211.t0 20.826
R16686 a_2672_211.n2 a_2672_211.n1 20.689
R16687 a_2577_196.n0 a_2577_196.t1 362.857
R16688 a_2577_196.t4 a_2577_196.t3 337.399
R16689 a_2577_196.t3 a_2577_196.t5 298.839
R16690 a_2577_196.n0 a_2577_196.t4 280.405
R16691 a_2577_196.n1 a_2577_196.t2 200
R16692 a_2577_196.n1 a_2577_196.n0 172.311
R16693 a_2577_196.n2 a_2577_196.n1 24
R16694 a_2577_196.n1 a_2577_196.t0 21.212
R16695 a_383_n953.n25 a_383_n953.t27 561.971
R16696 a_383_n953.n0 a_383_n953.t4 461.908
R16697 a_383_n953.t12 a_383_n953.n25 108.635
R16698 a_383_n953.n0 a_383_n953.t3 79.512
R16699 a_383_n953.n24 a_383_n953.t19 65.401
R16700 a_383_n953.n23 a_383_n953.t17 65.401
R16701 a_383_n953.n22 a_383_n953.t11 65.401
R16702 a_383_n953.n21 a_383_n953.t13 65.401
R16703 a_383_n953.n20 a_383_n953.t22 65.401
R16704 a_383_n953.n19 a_383_n953.t15 65.401
R16705 a_383_n953.n18 a_383_n953.t16 65.401
R16706 a_383_n953.n17 a_383_n953.t9 65.401
R16707 a_383_n953.n16 a_383_n953.t2 65.401
R16708 a_383_n953.n15 a_383_n953.t7 65.401
R16709 a_383_n953.n14 a_383_n953.t20 65.401
R16710 a_383_n953.n13 a_383_n953.t23 65.401
R16711 a_383_n953.n12 a_383_n953.t14 65.401
R16712 a_383_n953.n11 a_383_n953.t5 65.401
R16713 a_383_n953.n10 a_383_n953.t10 65.401
R16714 a_383_n953.n9 a_383_n953.t21 65.401
R16715 a_383_n953.n8 a_383_n953.t18 65.401
R16716 a_383_n953.n7 a_383_n953.t1 65.401
R16717 a_383_n953.n6 a_383_n953.t0 65.401
R16718 a_383_n953.n5 a_383_n953.t26 65.401
R16719 a_383_n953.n4 a_383_n953.t8 65.401
R16720 a_383_n953.n3 a_383_n953.t24 65.401
R16721 a_383_n953.n2 a_383_n953.t25 65.401
R16722 a_383_n953.n1 a_383_n953.t6 65.401
R16723 a_383_n953.n1 a_383_n953.n0 5.64
R16724 a_383_n953.n25 a_383_n953.n24 4.438
R16725 a_383_n953.n23 a_383_n953.n22 2.524
R16726 a_383_n953.n3 a_383_n953.n2 2.498
R16727 a_383_n953.n17 a_383_n953.n16 2.364
R16728 a_383_n953.n9 a_383_n953.n8 2.355
R16729 a_383_n953.n2 a_383_n953.n1 1.998
R16730 a_383_n953.n4 a_383_n953.n3 1.998
R16731 a_383_n953.n5 a_383_n953.n4 1.998
R16732 a_383_n953.n6 a_383_n953.n5 1.998
R16733 a_383_n953.n7 a_383_n953.n6 1.998
R16734 a_383_n953.n8 a_383_n953.n7 1.998
R16735 a_383_n953.n10 a_383_n953.n9 1.998
R16736 a_383_n953.n11 a_383_n953.n10 1.998
R16737 a_383_n953.n12 a_383_n953.n11 1.998
R16738 a_383_n953.n13 a_383_n953.n12 1.998
R16739 a_383_n953.n14 a_383_n953.n13 1.998
R16740 a_383_n953.n15 a_383_n953.n14 1.998
R16741 a_383_n953.n16 a_383_n953.n15 1.998
R16742 a_383_n953.n18 a_383_n953.n17 1.998
R16743 a_383_n953.n19 a_383_n953.n18 1.998
R16744 a_383_n953.n20 a_383_n953.n19 1.998
R16745 a_383_n953.n21 a_383_n953.n20 1.998
R16746 a_383_n953.n22 a_383_n953.n21 1.998
R16747 a_383_n953.n24 a_383_n953.n23 1.998
R16748 a_7306_n8026.t1 a_7306_n8026.t0 336.814
R16749 a_7247_n8071.t0 a_7247_n8071.t1 68.74
R16750 a_8221_n8583.n0 a_8221_n8583.t4 1465.51
R16751 a_8221_n8583.n0 a_8221_n8583.t3 712.44
R16752 a_8221_n8583.n1 a_8221_n8583.t2 375.067
R16753 a_8221_n8583.n1 a_8221_n8583.t0 272.668
R16754 a_8221_n8583.n2 a_8221_n8583.n0 143.764
R16755 a_8221_n8583.t1 a_8221_n8583.n2 78.193
R16756 a_8221_n8583.n2 a_8221_n8583.n1 4.517
R16757 a_3231_n4378.n3 a_3231_n4378.t3 475.39
R16758 a_3231_n4378.n3 a_3231_n4378.n2 419.907
R16759 a_3231_n4378.t4 a_3231_n4378.t6 228.696
R16760 a_3231_n4378.n2 a_3231_n4378.t1 185.704
R16761 a_3231_n4378.n0 a_3231_n4378.t4 126.761
R16762 a_3231_n4378.n1 a_3231_n4378.t5 126.284
R16763 a_3231_n4378.n1 a_3231_n4378.t0 126.284
R16764 a_3231_n4378.t2 a_3231_n4378.n3 124.375
R16765 a_3231_n4378.t0 a_3231_n4378.n0 115.122
R16766 a_3231_n4378.n0 a_3231_n4378.t7 111.229
R16767 a_3231_n4378.n2 a_3231_n4378.n1 8.764
R16768 WWLD[2].n0 WWLD[2].t14 262.032
R16769 WWLD[2].n29 WWLD[2].t17 260.715
R16770 WWLD[2].n27 WWLD[2].t20 260.715
R16771 WWLD[2].n25 WWLD[2].t2 260.715
R16772 WWLD[2].n23 WWLD[2].t28 260.715
R16773 WWLD[2].n21 WWLD[2].t8 260.715
R16774 WWLD[2].n19 WWLD[2].t25 260.715
R16775 WWLD[2].n17 WWLD[2].t16 260.715
R16776 WWLD[2].n15 WWLD[2].t31 260.715
R16777 WWLD[2].n13 WWLD[2].t21 260.715
R16778 WWLD[2].n11 WWLD[2].t29 260.715
R16779 WWLD[2].n9 WWLD[2].t18 260.715
R16780 WWLD[2].n7 WWLD[2].t0 260.715
R16781 WWLD[2].n5 WWLD[2].t26 260.715
R16782 WWLD[2].n3 WWLD[2].t9 260.715
R16783 WWLD[2].n1 WWLD[2].t22 260.715
R16784 WWLD[2].n30 WWLD[2].t1 259.254
R16785 WWLD[2].n28 WWLD[2].t7 259.254
R16786 WWLD[2].n26 WWLD[2].t19 259.254
R16787 WWLD[2].n24 WWLD[2].t3 259.254
R16788 WWLD[2].n22 WWLD[2].t27 259.254
R16789 WWLD[2].n20 WWLD[2].t10 259.254
R16790 WWLD[2].n18 WWLD[2].t23 259.254
R16791 WWLD[2].n16 WWLD[2].t5 259.254
R16792 WWLD[2].n14 WWLD[2].t30 259.254
R16793 WWLD[2].n12 WWLD[2].t13 259.254
R16794 WWLD[2].n10 WWLD[2].t4 259.254
R16795 WWLD[2].n8 WWLD[2].t11 259.254
R16796 WWLD[2].n6 WWLD[2].t12 259.254
R16797 WWLD[2].n4 WWLD[2].t15 259.254
R16798 WWLD[2].n2 WWLD[2].t6 259.254
R16799 WWLD[2].n0 WWLD[2].t24 259.254
R16800 WWLD[2] WWLD[2].n30 44.647
R16801 WWLD[2].n1 WWLD[2].n0 3.576
R16802 WWLD[2].n3 WWLD[2].n2 3.576
R16803 WWLD[2].n5 WWLD[2].n4 3.576
R16804 WWLD[2].n7 WWLD[2].n6 3.576
R16805 WWLD[2].n9 WWLD[2].n8 3.576
R16806 WWLD[2].n11 WWLD[2].n10 3.576
R16807 WWLD[2].n13 WWLD[2].n12 3.576
R16808 WWLD[2].n15 WWLD[2].n14 3.576
R16809 WWLD[2].n17 WWLD[2].n16 3.576
R16810 WWLD[2].n19 WWLD[2].n18 3.576
R16811 WWLD[2].n21 WWLD[2].n20 3.576
R16812 WWLD[2].n23 WWLD[2].n22 3.576
R16813 WWLD[2].n25 WWLD[2].n24 3.576
R16814 WWLD[2].n27 WWLD[2].n26 3.576
R16815 WWLD[2].n29 WWLD[2].n28 3.576
R16816 WWLD[2].n2 WWLD[2].n1 1.317
R16817 WWLD[2].n4 WWLD[2].n3 1.317
R16818 WWLD[2].n6 WWLD[2].n5 1.317
R16819 WWLD[2].n8 WWLD[2].n7 1.317
R16820 WWLD[2].n10 WWLD[2].n9 1.317
R16821 WWLD[2].n12 WWLD[2].n11 1.317
R16822 WWLD[2].n14 WWLD[2].n13 1.317
R16823 WWLD[2].n16 WWLD[2].n15 1.317
R16824 WWLD[2].n18 WWLD[2].n17 1.317
R16825 WWLD[2].n20 WWLD[2].n19 1.317
R16826 WWLD[2].n22 WWLD[2].n21 1.317
R16827 WWLD[2].n24 WWLD[2].n23 1.317
R16828 WWLD[2].n26 WWLD[2].n25 1.317
R16829 WWLD[2].n28 WWLD[2].n27 1.317
R16830 WWLD[2].n30 WWLD[2].n29 1.317
R16831 a_6870_4887.n25 a_6870_4887.t27 561.971
R16832 a_6870_4887.n0 a_6870_4887.t4 449.944
R16833 a_6870_4887.t13 a_6870_4887.n25 108.636
R16834 a_6870_4887.n0 a_6870_4887.t3 74.821
R16835 a_6870_4887.n24 a_6870_4887.t21 63.519
R16836 a_6870_4887.n23 a_6870_4887.t19 63.519
R16837 a_6870_4887.n22 a_6870_4887.t12 63.519
R16838 a_6870_4887.n21 a_6870_4887.t14 63.519
R16839 a_6870_4887.n20 a_6870_4887.t24 63.519
R16840 a_6870_4887.n19 a_6870_4887.t17 63.519
R16841 a_6870_4887.n18 a_6870_4887.t18 63.519
R16842 a_6870_4887.n17 a_6870_4887.t10 63.519
R16843 a_6870_4887.n16 a_6870_4887.t2 63.519
R16844 a_6870_4887.n15 a_6870_4887.t8 63.519
R16845 a_6870_4887.n14 a_6870_4887.t22 63.519
R16846 a_6870_4887.n13 a_6870_4887.t5 63.519
R16847 a_6870_4887.n12 a_6870_4887.t16 63.519
R16848 a_6870_4887.n11 a_6870_4887.t6 63.519
R16849 a_6870_4887.n10 a_6870_4887.t11 63.519
R16850 a_6870_4887.n9 a_6870_4887.t23 63.519
R16851 a_6870_4887.n8 a_6870_4887.t20 63.519
R16852 a_6870_4887.n7 a_6870_4887.t1 63.519
R16853 a_6870_4887.n6 a_6870_4887.t0 63.519
R16854 a_6870_4887.n5 a_6870_4887.t26 63.519
R16855 a_6870_4887.n4 a_6870_4887.t9 63.519
R16856 a_6870_4887.n3 a_6870_4887.t15 63.519
R16857 a_6870_4887.n2 a_6870_4887.t25 63.519
R16858 a_6870_4887.n1 a_6870_4887.t7 63.519
R16859 a_6870_4887.n1 a_6870_4887.n0 8.619
R16860 a_6870_4887.n25 a_6870_4887.n24 2.946
R16861 a_6870_4887.n23 a_6870_4887.n22 2.524
R16862 a_6870_4887.n3 a_6870_4887.n2 2.498
R16863 a_6870_4887.n17 a_6870_4887.n16 2.364
R16864 a_6870_4887.n9 a_6870_4887.n8 2.355
R16865 a_6870_4887.n24 a_6870_4887.n23 1.998
R16866 a_6870_4887.n22 a_6870_4887.n21 1.998
R16867 a_6870_4887.n21 a_6870_4887.n20 1.998
R16868 a_6870_4887.n20 a_6870_4887.n19 1.998
R16869 a_6870_4887.n19 a_6870_4887.n18 1.998
R16870 a_6870_4887.n18 a_6870_4887.n17 1.998
R16871 a_6870_4887.n16 a_6870_4887.n15 1.998
R16872 a_6870_4887.n15 a_6870_4887.n14 1.998
R16873 a_6870_4887.n14 a_6870_4887.n13 1.998
R16874 a_6870_4887.n13 a_6870_4887.n12 1.998
R16875 a_6870_4887.n12 a_6870_4887.n11 1.998
R16876 a_6870_4887.n11 a_6870_4887.n10 1.998
R16877 a_6870_4887.n10 a_6870_4887.n9 1.998
R16878 a_6870_4887.n8 a_6870_4887.n7 1.998
R16879 a_6870_4887.n7 a_6870_4887.n6 1.998
R16880 a_6870_4887.n6 a_6870_4887.n5 1.998
R16881 a_6870_4887.n5 a_6870_4887.n4 1.998
R16882 a_6870_4887.n4 a_6870_4887.n3 1.998
R16883 a_6870_4887.n2 a_6870_4887.n1 1.998
R16884 a_6602_4133.n0 a_6602_4133.t1 362.857
R16885 a_6602_4133.t3 a_6602_4133.t5 337.399
R16886 a_6602_4133.t5 a_6602_4133.t4 298.839
R16887 a_6602_4133.n0 a_6602_4133.t3 280.405
R16888 a_6602_4133.n1 a_6602_4133.t0 200
R16889 a_6602_4133.n1 a_6602_4133.n0 172.311
R16890 a_6602_4133.n2 a_6602_4133.n1 24
R16891 a_6602_4133.n1 a_6602_4133.t2 21.212
R16892 a_7067_2943.t0 a_7067_2943.t1 242.857
R16893 a_2002_4430.n0 a_2002_4430.t1 362.857
R16894 a_2002_4430.t3 a_2002_4430.t5 337.399
R16895 a_2002_4430.t5 a_2002_4430.t4 298.839
R16896 a_2002_4430.n0 a_2002_4430.t3 280.405
R16897 a_2002_4430.n1 a_2002_4430.t2 200
R16898 a_2002_4430.n1 a_2002_4430.n0 172.311
R16899 a_2002_4430.n2 a_2002_4430.n1 24
R16900 a_2002_4430.n1 a_2002_4430.t0 21.212
R16901 a_2097_4445.n0 a_2097_4445.t1 358.166
R16902 a_2097_4445.t5 a_2097_4445.t3 337.399
R16903 a_2097_4445.t3 a_2097_4445.t4 285.986
R16904 a_2097_4445.n0 a_2097_4445.t5 282.573
R16905 a_2097_4445.n1 a_2097_4445.t2 202.857
R16906 a_2097_4445.n1 a_2097_4445.n0 173.817
R16907 a_2097_4445.n1 a_2097_4445.t0 20.826
R16908 a_2097_4445.n2 a_2097_4445.n1 20.689
R16909 a_1440_3907.t0 a_1440_3907.t1 242.857
R16910 a_4972_2421.n0 a_4972_2421.t2 358.166
R16911 a_4972_2421.t4 a_4972_2421.t3 337.399
R16912 a_4972_2421.t3 a_4972_2421.t5 285.986
R16913 a_4972_2421.n0 a_4972_2421.t4 282.573
R16914 a_4972_2421.n1 a_4972_2421.t0 202.857
R16915 a_4972_2421.n1 a_4972_2421.n0 173.817
R16916 a_4972_2421.n1 a_4972_2421.t1 20.826
R16917 a_4972_2421.n2 a_4972_2421.n1 20.689
R16918 a_2672_4148.n0 a_2672_4148.t1 358.166
R16919 a_2672_4148.t3 a_2672_4148.t4 337.399
R16920 a_2672_4148.t4 a_2672_4148.t5 285.986
R16921 a_2672_4148.n0 a_2672_4148.t3 282.573
R16922 a_2672_4148.n1 a_2672_4148.t0 202.857
R16923 a_2672_4148.n1 a_2672_4148.n0 173.817
R16924 a_2672_4148.n1 a_2672_4148.t2 20.826
R16925 a_2672_4148.n2 a_2672_4148.n1 20.689
R16926 a_2577_4133.n0 a_2577_4133.t2 362.857
R16927 a_2577_4133.t3 a_2577_4133.t4 337.399
R16928 a_2577_4133.t4 a_2577_4133.t5 298.839
R16929 a_2577_4133.n0 a_2577_4133.t3 280.405
R16930 a_2577_4133.n1 a_2577_4133.t0 200
R16931 a_2577_4133.n1 a_2577_4133.n0 172.311
R16932 a_2577_4133.n2 a_2577_4133.n1 24
R16933 a_2577_4133.n1 a_2577_4133.t1 21.212
R16934 a_3822_2180.n0 a_3822_2180.t0 358.166
R16935 a_3822_2180.t3 a_3822_2180.t5 337.399
R16936 a_3822_2180.t5 a_3822_2180.t4 285.986
R16937 a_3822_2180.n0 a_3822_2180.t3 282.573
R16938 a_3822_2180.n1 a_3822_2180.t2 202.857
R16939 a_3822_2180.n1 a_3822_2180.n0 173.817
R16940 a_3822_2180.n1 a_3822_2180.t1 20.826
R16941 a_3822_2180.n2 a_3822_2180.n1 20.689
R16942 a_3727_2165.n0 a_3727_2165.t1 362.857
R16943 a_3727_2165.t3 a_3727_2165.t4 337.399
R16944 a_3727_2165.t4 a_3727_2165.t5 298.839
R16945 a_3727_2165.n0 a_3727_2165.t3 280.405
R16946 a_3727_2165.n1 a_3727_2165.t2 200
R16947 a_3727_2165.n1 a_3727_2165.n0 172.311
R16948 a_3727_2165.n2 a_3727_2165.n1 24
R16949 a_3727_2165.n1 a_3727_2165.t0 21.212
R16950 a_4972_1939.n0 a_4972_1939.t2 358.166
R16951 a_4972_1939.t5 a_4972_1939.t4 337.399
R16952 a_4972_1939.t4 a_4972_1939.t3 285.986
R16953 a_4972_1939.n0 a_4972_1939.t5 282.573
R16954 a_4972_1939.n1 a_4972_1939.t0 202.857
R16955 a_4972_1939.n1 a_4972_1939.n0 173.817
R16956 a_4972_1939.n1 a_4972_1939.t1 20.826
R16957 a_4972_1939.n2 a_4972_1939.n1 20.689
R16958 a_372_452.n0 a_372_452.t0 358.166
R16959 a_372_452.t5 a_372_452.t4 337.399
R16960 a_372_452.t4 a_372_452.t3 285.986
R16961 a_372_452.n0 a_372_452.t5 282.573
R16962 a_372_452.n1 a_372_452.t2 202.857
R16963 a_372_452.n1 a_372_452.n0 173.817
R16964 a_372_452.n1 a_372_452.t1 20.826
R16965 a_372_452.n2 a_372_452.n1 20.689
R16966 a_742_452.t0 a_742_452.t1 242.857
R16967 a_13637_n3770.n0 a_13637_n3770.t0 65.064
R16968 a_13637_n3770.n0 a_13637_n3770.t2 42.011
R16969 a_13637_n3770.t1 a_13637_n3770.n0 2.113
R16970 a_4302_3410.n0 a_4302_3410.t1 362.857
R16971 a_4302_3410.t4 a_4302_3410.t3 337.399
R16972 a_4302_3410.t3 a_4302_3410.t5 298.839
R16973 a_4302_3410.n0 a_4302_3410.t4 280.405
R16974 a_4302_3410.n1 a_4302_3410.t0 200
R16975 a_4302_3410.n1 a_4302_3410.n0 172.311
R16976 a_4302_3410.n2 a_4302_3410.n1 24
R16977 a_4302_3410.n1 a_4302_3410.t2 21.212
R16978 a_4397_3425.n0 a_4397_3425.t2 358.166
R16979 a_4397_3425.t4 a_4397_3425.t5 337.399
R16980 a_4397_3425.t5 a_4397_3425.t3 285.986
R16981 a_4397_3425.n0 a_4397_3425.t4 282.573
R16982 a_4397_3425.n1 a_4397_3425.t0 202.857
R16983 a_4397_3425.n1 a_4397_3425.n0 173.817
R16984 a_4397_3425.n1 a_4397_3425.t1 20.826
R16985 a_4397_3425.n2 a_4397_3425.n1 20.689
R16986 a_8410_n1770.n0 a_8410_n1770.t1 325.682
R16987 a_8410_n1770.n0 a_8410_n1770.t2 322.294
R16988 a_8410_n1770.t0 a_8410_n1770.n0 73.623
R16989 a_8452_n1770.t0 a_8452_n1770.t1 213.924
R16990 a_2590_n1053.t0 a_2590_n1053.t1 242.857
R16991 a_3247_452.n0 a_3247_452.t2 358.166
R16992 a_3247_452.t3 a_3247_452.t5 337.399
R16993 a_3247_452.t5 a_3247_452.t4 285.986
R16994 a_3247_452.n0 a_3247_452.t3 282.573
R16995 a_3247_452.n1 a_3247_452.t0 202.857
R16996 a_3247_452.n1 a_3247_452.n0 173.817
R16997 a_3247_452.n1 a_3247_452.t1 20.826
R16998 a_3247_452.n2 a_3247_452.n1 20.689
R16999 a_3152_437.n0 a_3152_437.t1 362.857
R17000 a_3152_437.t4 a_3152_437.t3 337.399
R17001 a_3152_437.t3 a_3152_437.t5 298.839
R17002 a_3152_437.n0 a_3152_437.t4 280.405
R17003 a_3152_437.n1 a_3152_437.t2 200
R17004 a_3152_437.n1 a_3152_437.n0 172.311
R17005 a_3152_437.n2 a_3152_437.n1 24
R17006 a_3152_437.n1 a_3152_437.t0 21.212
R17007 ADC0_OUT[2].n0 ADC0_OUT[2].t4 1354.27
R17008 ADC0_OUT[2].n0 ADC0_OUT[2].t3 821.954
R17009 ADC0_OUT[2].n3 ADC0_OUT[2].t0 349.397
R17010 ADC0_OUT[2].n2 ADC0_OUT[2].t1 266.575
R17011 ADC0_OUT[2].n1 ADC0_OUT[2].n0 149.035
R17012 ADC0_OUT[2].n1 ADC0_OUT[2].t2 46.723
R17013 ADC0_OUT[2] ADC0_OUT[2].n3 38.04
R17014 ADC0_OUT[2].n3 ADC0_OUT[2].n2 34.635
R17015 ADC0_OUT[2].n2 ADC0_OUT[2].n1 17.317
R17016 RWLB[10].n0 RWLB[10].t13 154.228
R17017 RWLB[10].n14 RWLB[10].t14 149.249
R17018 RWLB[10].n13 RWLB[10].t0 149.249
R17019 RWLB[10].n12 RWLB[10].t11 149.249
R17020 RWLB[10].n11 RWLB[10].t5 149.249
R17021 RWLB[10].n10 RWLB[10].t15 149.249
R17022 RWLB[10].n9 RWLB[10].t2 149.249
R17023 RWLB[10].n8 RWLB[10].t3 149.249
R17024 RWLB[10].n7 RWLB[10].t8 149.249
R17025 RWLB[10].n6 RWLB[10].t1 149.249
R17026 RWLB[10].n5 RWLB[10].t6 149.249
R17027 RWLB[10].n4 RWLB[10].t7 149.249
R17028 RWLB[10].n3 RWLB[10].t12 149.249
R17029 RWLB[10].n2 RWLB[10].t4 149.249
R17030 RWLB[10].n1 RWLB[10].t10 149.249
R17031 RWLB[10].n0 RWLB[10].t9 149.249
R17032 RWLB[10] RWLB[10].n14 47.816
R17033 RWLB[10].n1 RWLB[10].n0 4.979
R17034 RWLB[10].n2 RWLB[10].n1 4.979
R17035 RWLB[10].n3 RWLB[10].n2 4.979
R17036 RWLB[10].n4 RWLB[10].n3 4.979
R17037 RWLB[10].n5 RWLB[10].n4 4.979
R17038 RWLB[10].n6 RWLB[10].n5 4.979
R17039 RWLB[10].n7 RWLB[10].n6 4.979
R17040 RWLB[10].n8 RWLB[10].n7 4.979
R17041 RWLB[10].n9 RWLB[10].n8 4.979
R17042 RWLB[10].n10 RWLB[10].n9 4.979
R17043 RWLB[10].n11 RWLB[10].n10 4.979
R17044 RWLB[10].n12 RWLB[10].n11 4.979
R17045 RWLB[10].n13 RWLB[10].n12 4.979
R17046 RWLB[10].n14 RWLB[10].n13 4.979
R17047 a_1317_1216.t0 a_1317_1216.t1 242.857
R17048 WWLD[6].n0 WWLD[6].t28 262.032
R17049 WWLD[6].n29 WWLD[6].t31 260.715
R17050 WWLD[6].n27 WWLD[6].t1 260.715
R17051 WWLD[6].n25 WWLD[6].t21 260.715
R17052 WWLD[6].n23 WWLD[6].t12 260.715
R17053 WWLD[6].n21 WWLD[6].t23 260.715
R17054 WWLD[6].n19 WWLD[6].t7 260.715
R17055 WWLD[6].n17 WWLD[6].t30 260.715
R17056 WWLD[6].n15 WWLD[6].t17 260.715
R17057 WWLD[6].n13 WWLD[6].t3 260.715
R17058 WWLD[6].n11 WWLD[6].t13 260.715
R17059 WWLD[6].n9 WWLD[6].t0 260.715
R17060 WWLD[6].n7 WWLD[6].t19 260.715
R17061 WWLD[6].n5 WWLD[6].t8 260.715
R17062 WWLD[6].n3 WWLD[6].t24 260.715
R17063 WWLD[6].n1 WWLD[6].t4 260.715
R17064 WWLD[6].n30 WWLD[6].t2 259.254
R17065 WWLD[6].n28 WWLD[6].t11 259.254
R17066 WWLD[6].n26 WWLD[6].t22 259.254
R17067 WWLD[6].n24 WWLD[6].t5 259.254
R17068 WWLD[6].n22 WWLD[6].t27 259.254
R17069 WWLD[6].n20 WWLD[6].t14 259.254
R17070 WWLD[6].n18 WWLD[6].t25 259.254
R17071 WWLD[6].n16 WWLD[6].t9 259.254
R17072 WWLD[6].n14 WWLD[6].t29 259.254
R17073 WWLD[6].n12 WWLD[6].t18 259.254
R17074 WWLD[6].n10 WWLD[6].t6 259.254
R17075 WWLD[6].n8 WWLD[6].t15 259.254
R17076 WWLD[6].n6 WWLD[6].t16 259.254
R17077 WWLD[6].n4 WWLD[6].t20 259.254
R17078 WWLD[6].n2 WWLD[6].t10 259.254
R17079 WWLD[6].n0 WWLD[6].t26 259.254
R17080 WWLD[6] WWLD[6].n30 44.647
R17081 WWLD[6].n1 WWLD[6].n0 3.576
R17082 WWLD[6].n3 WWLD[6].n2 3.576
R17083 WWLD[6].n5 WWLD[6].n4 3.576
R17084 WWLD[6].n7 WWLD[6].n6 3.576
R17085 WWLD[6].n9 WWLD[6].n8 3.576
R17086 WWLD[6].n11 WWLD[6].n10 3.576
R17087 WWLD[6].n13 WWLD[6].n12 3.576
R17088 WWLD[6].n15 WWLD[6].n14 3.576
R17089 WWLD[6].n17 WWLD[6].n16 3.576
R17090 WWLD[6].n19 WWLD[6].n18 3.576
R17091 WWLD[6].n21 WWLD[6].n20 3.576
R17092 WWLD[6].n23 WWLD[6].n22 3.576
R17093 WWLD[6].n25 WWLD[6].n24 3.576
R17094 WWLD[6].n27 WWLD[6].n26 3.576
R17095 WWLD[6].n29 WWLD[6].n28 3.576
R17096 WWLD[6].n2 WWLD[6].n1 1.317
R17097 WWLD[6].n4 WWLD[6].n3 1.317
R17098 WWLD[6].n6 WWLD[6].n5 1.317
R17099 WWLD[6].n8 WWLD[6].n7 1.317
R17100 WWLD[6].n10 WWLD[6].n9 1.317
R17101 WWLD[6].n12 WWLD[6].n11 1.317
R17102 WWLD[6].n14 WWLD[6].n13 1.317
R17103 WWLD[6].n16 WWLD[6].n15 1.317
R17104 WWLD[6].n18 WWLD[6].n17 1.317
R17105 WWLD[6].n20 WWLD[6].n19 1.317
R17106 WWLD[6].n22 WWLD[6].n21 1.317
R17107 WWLD[6].n24 WWLD[6].n23 1.317
R17108 WWLD[6].n26 WWLD[6].n25 1.317
R17109 WWLD[6].n28 WWLD[6].n27 1.317
R17110 WWLD[6].n30 WWLD[6].n29 1.317
R17111 a_6295_4887.n25 a_6295_4887.t27 561.971
R17112 a_6295_4887.n0 a_6295_4887.t5 449.944
R17113 a_6295_4887.t12 a_6295_4887.n25 108.636
R17114 a_6295_4887.n0 a_6295_4887.t4 74.821
R17115 a_6295_4887.n24 a_6295_4887.t19 63.519
R17116 a_6295_4887.n23 a_6295_4887.t0 63.519
R17117 a_6295_4887.n22 a_6295_4887.t11 63.519
R17118 a_6295_4887.n21 a_6295_4887.t13 63.519
R17119 a_6295_4887.n20 a_6295_4887.t24 63.519
R17120 a_6295_4887.n19 a_6295_4887.t16 63.519
R17121 a_6295_4887.n18 a_6295_4887.t17 63.519
R17122 a_6295_4887.n17 a_6295_4887.t9 63.519
R17123 a_6295_4887.n16 a_6295_4887.t3 63.519
R17124 a_6295_4887.n15 a_6295_4887.t7 63.519
R17125 a_6295_4887.n14 a_6295_4887.t20 63.519
R17126 a_6295_4887.n13 a_6295_4887.t22 63.519
R17127 a_6295_4887.n12 a_6295_4887.t15 63.519
R17128 a_6295_4887.n11 a_6295_4887.t25 63.519
R17129 a_6295_4887.n10 a_6295_4887.t10 63.519
R17130 a_6295_4887.n9 a_6295_4887.t21 63.519
R17131 a_6295_4887.n8 a_6295_4887.t18 63.519
R17132 a_6295_4887.n7 a_6295_4887.t2 63.519
R17133 a_6295_4887.n6 a_6295_4887.t1 63.519
R17134 a_6295_4887.n5 a_6295_4887.t26 63.519
R17135 a_6295_4887.n4 a_6295_4887.t8 63.519
R17136 a_6295_4887.n3 a_6295_4887.t14 63.519
R17137 a_6295_4887.n2 a_6295_4887.t23 63.519
R17138 a_6295_4887.n1 a_6295_4887.t6 63.519
R17139 a_6295_4887.n1 a_6295_4887.n0 8.619
R17140 a_6295_4887.n25 a_6295_4887.n24 2.946
R17141 a_6295_4887.n23 a_6295_4887.n22 2.524
R17142 a_6295_4887.n3 a_6295_4887.n2 2.498
R17143 a_6295_4887.n17 a_6295_4887.n16 2.364
R17144 a_6295_4887.n9 a_6295_4887.n8 2.355
R17145 a_6295_4887.n24 a_6295_4887.n23 1.998
R17146 a_6295_4887.n22 a_6295_4887.n21 1.998
R17147 a_6295_4887.n21 a_6295_4887.n20 1.998
R17148 a_6295_4887.n20 a_6295_4887.n19 1.998
R17149 a_6295_4887.n19 a_6295_4887.n18 1.998
R17150 a_6295_4887.n18 a_6295_4887.n17 1.998
R17151 a_6295_4887.n16 a_6295_4887.n15 1.998
R17152 a_6295_4887.n15 a_6295_4887.n14 1.998
R17153 a_6295_4887.n14 a_6295_4887.n13 1.998
R17154 a_6295_4887.n13 a_6295_4887.n12 1.998
R17155 a_6295_4887.n12 a_6295_4887.n11 1.998
R17156 a_6295_4887.n11 a_6295_4887.n10 1.998
R17157 a_6295_4887.n10 a_6295_4887.n9 1.998
R17158 a_6295_4887.n8 a_6295_4887.n7 1.998
R17159 a_6295_4887.n7 a_6295_4887.n6 1.998
R17160 a_6295_4887.n6 a_6295_4887.n5 1.998
R17161 a_6295_4887.n5 a_6295_4887.n4 1.998
R17162 a_6295_4887.n4 a_6295_4887.n3 1.998
R17163 a_6295_4887.n2 a_6295_4887.n1 1.998
R17164 a_6027_n827.n0 a_6027_n827.t2 362.857
R17165 a_6027_n827.t3 a_6027_n827.t4 337.399
R17166 a_6027_n827.t4 a_6027_n827.t5 298.839
R17167 a_6027_n827.n0 a_6027_n827.t3 280.405
R17168 a_6027_n827.n1 a_6027_n827.t0 200
R17169 a_6027_n827.n1 a_6027_n827.n0 172.311
R17170 a_6027_n827.n2 a_6027_n827.n1 24
R17171 a_6027_n827.n1 a_6027_n827.t1 21.212
R17172 a_8902_196.n0 a_8902_196.t2 362.857
R17173 a_8902_196.t5 a_8902_196.t4 337.399
R17174 a_8902_196.t4 a_8902_196.t3 298.839
R17175 a_8902_196.n0 a_8902_196.t5 280.405
R17176 a_8902_196.n1 a_8902_196.t1 200
R17177 a_8902_196.n1 a_8902_196.n0 172.311
R17178 a_8902_196.n2 a_8902_196.n1 24
R17179 a_8902_196.n1 a_8902_196.t0 21.212
R17180 a_n3565_n5850.n0 a_n3565_n5850.t4 1465.51
R17181 a_n3565_n5850.n0 a_n3565_n5850.t3 712.44
R17182 a_n3565_n5850.n1 a_n3565_n5850.t0 375.067
R17183 a_n3565_n5850.n1 a_n3565_n5850.t1 272.668
R17184 a_n3565_n5850.n2 a_n3565_n5850.n0 143.764
R17185 a_n3565_n5850.t2 a_n3565_n5850.n2 78.193
R17186 a_n3565_n5850.n2 a_n3565_n5850.n1 4.517
R17187 a_11549_n3770.n0 a_11549_n3770.t0 65.064
R17188 a_11549_n3770.t1 a_11549_n3770.n0 42.011
R17189 a_11549_n3770.n0 a_11549_n3770.t2 2.113
R17190 a_8422_2180.n0 a_8422_2180.t1 358.166
R17191 a_8422_2180.t4 a_8422_2180.t3 337.399
R17192 a_8422_2180.t3 a_8422_2180.t5 285.986
R17193 a_8422_2180.n0 a_8422_2180.t4 282.573
R17194 a_8422_2180.n1 a_8422_2180.t2 202.857
R17195 a_8422_2180.n1 a_8422_2180.n0 173.817
R17196 a_8422_2180.n1 a_8422_2180.t0 20.826
R17197 a_8422_2180.n2 a_8422_2180.n1 20.689
R17198 a_8327_2165.n0 a_8327_2165.t1 362.857
R17199 a_8327_2165.t4 a_8327_2165.t5 337.399
R17200 a_8327_2165.t5 a_8327_2165.t3 298.839
R17201 a_8327_2165.n0 a_8327_2165.t4 280.405
R17202 a_8327_2165.n1 a_8327_2165.t2 200
R17203 a_8327_2165.n1 a_8327_2165.n0 172.311
R17204 a_8327_2165.n2 a_8327_2165.n1 24
R17205 a_8327_2165.n1 a_8327_2165.t0 21.212
R17206 RWL[8].n0 RWL[8].t4 154.243
R17207 RWL[8].n14 RWL[8].t10 149.249
R17208 RWL[8].n13 RWL[8].t15 149.249
R17209 RWL[8].n12 RWL[8].t6 149.249
R17210 RWL[8].n11 RWL[8].t11 149.249
R17211 RWL[8].n10 RWL[8].t8 149.249
R17212 RWL[8].n9 RWL[8].t0 149.249
R17213 RWL[8].n8 RWL[8].t7 149.249
R17214 RWL[8].n7 RWL[8].t13 149.249
R17215 RWL[8].n6 RWL[8].t9 149.249
R17216 RWL[8].n5 RWL[8].t3 149.249
R17217 RWL[8].n4 RWL[8].t12 149.249
R17218 RWL[8].n3 RWL[8].t1 149.249
R17219 RWL[8].n2 RWL[8].t2 149.249
R17220 RWL[8].n1 RWL[8].t5 149.249
R17221 RWL[8].n0 RWL[8].t14 149.249
R17222 RWL[8] RWL[8].n14 42.872
R17223 RWL[8].n1 RWL[8].n0 4.994
R17224 RWL[8].n2 RWL[8].n1 4.994
R17225 RWL[8].n3 RWL[8].n2 4.994
R17226 RWL[8].n4 RWL[8].n3 4.994
R17227 RWL[8].n5 RWL[8].n4 4.994
R17228 RWL[8].n6 RWL[8].n5 4.994
R17229 RWL[8].n7 RWL[8].n6 4.994
R17230 RWL[8].n8 RWL[8].n7 4.994
R17231 RWL[8].n9 RWL[8].n8 4.994
R17232 RWL[8].n10 RWL[8].n9 4.994
R17233 RWL[8].n11 RWL[8].n10 4.994
R17234 RWL[8].n12 RWL[8].n11 4.994
R17235 RWL[8].n13 RWL[8].n12 4.994
R17236 RWL[8].n14 RWL[8].n13 4.994
R17237 a_3165_1698.t0 a_3165_1698.t1 242.857
R17238 a_6027_1683.n0 a_6027_1683.t1 362.857
R17239 a_6027_1683.t5 a_6027_1683.t3 337.399
R17240 a_6027_1683.t3 a_6027_1683.t4 298.839
R17241 a_6027_1683.n0 a_6027_1683.t5 280.405
R17242 a_6027_1683.n1 a_6027_1683.t2 200
R17243 a_6027_1683.n1 a_6027_1683.n0 172.311
R17244 a_6027_1683.n2 a_6027_1683.n1 24
R17245 a_6027_1683.n1 a_6027_1683.t0 21.212
R17246 a_6122_1698.n0 a_6122_1698.t2 358.166
R17247 a_6122_1698.t4 a_6122_1698.t3 337.399
R17248 a_6122_1698.t3 a_6122_1698.t5 285.986
R17249 a_6122_1698.n0 a_6122_1698.t4 282.573
R17250 a_6122_1698.n1 a_6122_1698.t0 202.857
R17251 a_6122_1698.n1 a_6122_1698.n0 173.817
R17252 a_6122_1698.n1 a_6122_1698.t1 20.826
R17253 a_6122_1698.n2 a_6122_1698.n1 20.689
R17254 a_277_n45.n0 a_277_n45.t0 362.857
R17255 a_277_n45.t5 a_277_n45.t4 337.399
R17256 a_277_n45.t4 a_277_n45.t3 298.839
R17257 a_277_n45.n0 a_277_n45.t5 280.405
R17258 a_277_n45.n1 a_277_n45.t1 200
R17259 a_277_n45.n1 a_277_n45.n0 172.311
R17260 a_277_n45.n2 a_277_n45.n1 24
R17261 a_277_n45.n1 a_277_n45.t2 21.212
R17262 a_290_n30.t0 a_290_n30.t1 242.857
R17263 a_6693_n2422.n3 a_6693_n2422.t3 475.39
R17264 a_6693_n2422.n3 a_6693_n2422.n2 318.091
R17265 a_6693_n2422.t4 a_6693_n2422.t6 228.696
R17266 a_6693_n2422.n2 a_6693_n2422.t1 185.704
R17267 a_6693_n2422.n0 a_6693_n2422.t4 126.761
R17268 a_6693_n2422.n1 a_6693_n2422.t5 126.284
R17269 a_6693_n2422.n1 a_6693_n2422.t0 126.284
R17270 a_6693_n2422.t2 a_6693_n2422.n3 124.375
R17271 a_6693_n2422.t0 a_6693_n2422.n0 115.122
R17272 a_6693_n2422.n0 a_6693_n2422.t7 111.229
R17273 a_6693_n2422.n2 a_6693_n2422.n1 8.764
R17274 a_7272_4148.n0 a_7272_4148.t2 358.166
R17275 a_7272_4148.t4 a_7272_4148.t3 337.399
R17276 a_7272_4148.t3 a_7272_4148.t5 285.986
R17277 a_7272_4148.n0 a_7272_4148.t4 282.573
R17278 a_7272_4148.n1 a_7272_4148.t0 202.857
R17279 a_7272_4148.n1 a_7272_4148.n0 173.817
R17280 a_7272_4148.n1 a_7272_4148.t1 20.826
R17281 a_7272_4148.n2 a_7272_4148.n1 20.689
R17282 a_7177_4133.n0 a_7177_4133.t1 362.857
R17283 a_7177_4133.t5 a_7177_4133.t3 337.399
R17284 a_7177_4133.t3 a_7177_4133.t4 298.839
R17285 a_7177_4133.n0 a_7177_4133.t5 280.405
R17286 a_7177_4133.n1 a_7177_4133.t2 200
R17287 a_7177_4133.n1 a_7177_4133.n0 172.311
R17288 a_7177_4133.n2 a_7177_4133.n1 24
R17289 a_7177_4133.n1 a_7177_4133.t0 21.212
R17290 a_2015_3666.t0 a_2015_3666.t1 242.857
R17291 a_1317_211.t0 a_1317_211.t1 242.857
R17292 a_n3495_n4470.n0 a_n3495_n4470.t0 63.08
R17293 a_n3495_n4470.n0 a_n3495_n4470.t2 41.305
R17294 a_n3495_n4470.t1 a_n3495_n4470.n0 2.251
R17295 a_n3357_n4470.t0 a_n3357_n4470.t1 68.741
R17296 a_4972_3184.n0 a_4972_3184.t2 358.166
R17297 a_4972_3184.t4 a_4972_3184.t3 337.399
R17298 a_4972_3184.t3 a_4972_3184.t5 285.986
R17299 a_4972_3184.n0 a_4972_3184.t4 282.573
R17300 a_4972_3184.n1 a_4972_3184.t1 202.857
R17301 a_4972_3184.n1 a_4972_3184.n0 173.817
R17302 a_4972_3184.n1 a_4972_3184.t0 20.826
R17303 a_4972_3184.n2 a_4972_3184.n1 20.689
R17304 a_4983_n953.n25 a_4983_n953.t27 561.971
R17305 a_4983_n953.n0 a_4983_n953.t5 461.908
R17306 a_4983_n953.t13 a_4983_n953.n25 108.635
R17307 a_4983_n953.n0 a_4983_n953.t6 79.512
R17308 a_4983_n953.n24 a_4983_n953.t20 65.401
R17309 a_4983_n953.n23 a_4983_n953.t0 65.401
R17310 a_4983_n953.n22 a_4983_n953.t12 65.401
R17311 a_4983_n953.n21 a_4983_n953.t14 65.401
R17312 a_4983_n953.n20 a_4983_n953.t24 65.401
R17313 a_4983_n953.n19 a_4983_n953.t17 65.401
R17314 a_4983_n953.n18 a_4983_n953.t18 65.401
R17315 a_4983_n953.n17 a_4983_n953.t10 65.401
R17316 a_4983_n953.n16 a_4983_n953.t4 65.401
R17317 a_4983_n953.n15 a_4983_n953.t8 65.401
R17318 a_4983_n953.n14 a_4983_n953.t21 65.401
R17319 a_4983_n953.n13 a_4983_n953.t1 65.401
R17320 a_4983_n953.n12 a_4983_n953.t16 65.401
R17321 a_4983_n953.n11 a_4983_n953.t25 65.401
R17322 a_4983_n953.n10 a_4983_n953.t11 65.401
R17323 a_4983_n953.n9 a_4983_n953.t22 65.401
R17324 a_4983_n953.n8 a_4983_n953.t19 65.401
R17325 a_4983_n953.n7 a_4983_n953.t3 65.401
R17326 a_4983_n953.n6 a_4983_n953.t2 65.401
R17327 a_4983_n953.n5 a_4983_n953.t26 65.401
R17328 a_4983_n953.n4 a_4983_n953.t9 65.401
R17329 a_4983_n953.n3 a_4983_n953.t15 65.401
R17330 a_4983_n953.n2 a_4983_n953.t23 65.401
R17331 a_4983_n953.n1 a_4983_n953.t7 65.401
R17332 a_4983_n953.n1 a_4983_n953.n0 5.64
R17333 a_4983_n953.n25 a_4983_n953.n24 4.438
R17334 a_4983_n953.n23 a_4983_n953.n22 2.524
R17335 a_4983_n953.n3 a_4983_n953.n2 2.498
R17336 a_4983_n953.n17 a_4983_n953.n16 2.364
R17337 a_4983_n953.n9 a_4983_n953.n8 2.355
R17338 a_4983_n953.n2 a_4983_n953.n1 1.998
R17339 a_4983_n953.n4 a_4983_n953.n3 1.998
R17340 a_4983_n953.n5 a_4983_n953.n4 1.998
R17341 a_4983_n953.n6 a_4983_n953.n5 1.998
R17342 a_4983_n953.n7 a_4983_n953.n6 1.998
R17343 a_4983_n953.n8 a_4983_n953.n7 1.998
R17344 a_4983_n953.n10 a_4983_n953.n9 1.998
R17345 a_4983_n953.n11 a_4983_n953.n10 1.998
R17346 a_4983_n953.n12 a_4983_n953.n11 1.998
R17347 a_4983_n953.n13 a_4983_n953.n12 1.998
R17348 a_4983_n953.n14 a_4983_n953.n13 1.998
R17349 a_4983_n953.n15 a_4983_n953.n14 1.998
R17350 a_4983_n953.n16 a_4983_n953.n15 1.998
R17351 a_4983_n953.n18 a_4983_n953.n17 1.998
R17352 a_4983_n953.n19 a_4983_n953.n18 1.998
R17353 a_4983_n953.n20 a_4983_n953.n19 1.998
R17354 a_4983_n953.n21 a_4983_n953.n20 1.998
R17355 a_4983_n953.n22 a_4983_n953.n21 1.998
R17356 a_4983_n953.n24 a_4983_n953.n23 1.998
R17357 a_2381_n5338.n0 a_2381_n5338.t0 63.08
R17358 a_2381_n5338.n0 a_2381_n5338.t2 41.307
R17359 a_2381_n5338.t1 a_2381_n5338.n0 2.251
R17360 a_2519_n5338.t0 a_2519_n5338.t1 68.74
R17361 a_7177_3410.n0 a_7177_3410.t2 362.857
R17362 a_7177_3410.t4 a_7177_3410.t5 337.399
R17363 a_7177_3410.t5 a_7177_3410.t3 298.839
R17364 a_7177_3410.n0 a_7177_3410.t4 280.405
R17365 a_7177_3410.n1 a_7177_3410.t0 200
R17366 a_7177_3410.n1 a_7177_3410.n0 172.311
R17367 a_7177_3410.n2 a_7177_3410.n1 24
R17368 a_7177_3410.n1 a_7177_3410.t1 21.212
R17369 a_7190_3425.t0 a_7190_3425.t1 242.857
R17370 a_852_1924.n0 a_852_1924.t1 362.857
R17371 a_852_1924.t3 a_852_1924.t4 337.399
R17372 a_852_1924.t4 a_852_1924.t5 298.839
R17373 a_852_1924.n0 a_852_1924.t3 280.405
R17374 a_852_1924.n1 a_852_1924.t2 200
R17375 a_852_1924.n1 a_852_1924.n0 172.311
R17376 a_852_1924.n2 a_852_1924.n1 24
R17377 a_852_1924.n1 a_852_1924.t0 21.212
R17378 a_8902_437.n0 a_8902_437.t0 362.857
R17379 a_8902_437.t3 a_8902_437.t5 337.399
R17380 a_8902_437.t5 a_8902_437.t4 298.839
R17381 a_8902_437.n0 a_8902_437.t3 280.405
R17382 a_8902_437.n1 a_8902_437.t2 200
R17383 a_8902_437.n1 a_8902_437.n0 172.311
R17384 a_8902_437.n2 a_8902_437.n1 24
R17385 a_8902_437.n1 a_8902_437.t1 21.212
R17386 a_8997_452.n0 a_8997_452.t2 358.166
R17387 a_8997_452.t4 a_8997_452.t3 337.399
R17388 a_8997_452.t3 a_8997_452.t5 285.986
R17389 a_8997_452.n0 a_8997_452.t4 282.573
R17390 a_8997_452.n1 a_8997_452.t0 202.857
R17391 a_8997_452.n1 a_8997_452.n0 173.817
R17392 a_8997_452.n1 a_8997_452.t1 20.826
R17393 a_8997_452.n2 a_8997_452.n1 20.689
R17394 a_3165_n812.t0 a_3165_n812.t1 242.857
R17395 a_5118_n2426.n3 a_5118_n2426.n2 480.868
R17396 a_5118_n2426.n3 a_5118_n2426.t3 475.39
R17397 a_5118_n2426.t5 a_5118_n2426.t7 228.696
R17398 a_5118_n2426.n2 a_5118_n2426.t1 185.704
R17399 a_5118_n2426.n0 a_5118_n2426.t5 126.761
R17400 a_5118_n2426.n1 a_5118_n2426.t6 126.284
R17401 a_5118_n2426.n1 a_5118_n2426.t0 126.284
R17402 a_5118_n2426.t2 a_5118_n2426.n3 124.375
R17403 a_5118_n2426.t0 a_5118_n2426.n0 115.122
R17404 a_5118_n2426.n0 a_5118_n2426.t4 111.229
R17405 a_5118_n2426.n2 a_5118_n2426.n1 8.764
R17406 a_5595_n5092.t0 a_5595_n5092.t1 42.705
R17407 a_n1163_n4470.n0 a_n1163_n4470.t0 63.08
R17408 a_n1163_n4470.n0 a_n1163_n4470.t2 41.305
R17409 a_n1163_n4470.t1 a_n1163_n4470.n0 2.251
R17410 WWL[4].n0 WWL[4].t0 262.032
R17411 WWL[4].n29 WWL[4].t3 260.715
R17412 WWL[4].n27 WWL[4].t6 260.715
R17413 WWL[4].n25 WWL[4].t20 260.715
R17414 WWL[4].n23 WWL[4].t14 260.715
R17415 WWL[4].n21 WWL[4].t26 260.715
R17416 WWL[4].n19 WWL[4].t11 260.715
R17417 WWL[4].n17 WWL[4].t2 260.715
R17418 WWL[4].n15 WWL[4].t17 260.715
R17419 WWL[4].n13 WWL[4].t7 260.715
R17420 WWL[4].n11 WWL[4].t15 260.715
R17421 WWL[4].n9 WWL[4].t4 260.715
R17422 WWL[4].n7 WWL[4].t18 260.715
R17423 WWL[4].n5 WWL[4].t12 260.715
R17424 WWL[4].n3 WWL[4].t27 260.715
R17425 WWL[4].n1 WWL[4].t8 260.715
R17426 WWL[4].n30 WWL[4].t19 259.254
R17427 WWL[4].n28 WWL[4].t25 259.254
R17428 WWL[4].n26 WWL[4].t5 259.254
R17429 WWL[4].n24 WWL[4].t21 259.254
R17430 WWL[4].n22 WWL[4].t13 259.254
R17431 WWL[4].n20 WWL[4].t28 259.254
R17432 WWL[4].n18 WWL[4].t9 259.254
R17433 WWL[4].n16 WWL[4].t23 259.254
R17434 WWL[4].n14 WWL[4].t16 259.254
R17435 WWL[4].n12 WWL[4].t31 259.254
R17436 WWL[4].n10 WWL[4].t22 259.254
R17437 WWL[4].n8 WWL[4].t29 259.254
R17438 WWL[4].n6 WWL[4].t30 259.254
R17439 WWL[4].n4 WWL[4].t1 259.254
R17440 WWL[4].n2 WWL[4].t24 259.254
R17441 WWL[4].n0 WWL[4].t10 259.254
R17442 WWL[4] WWL[4].n30 44.647
R17443 WWL[4].n1 WWL[4].n0 3.576
R17444 WWL[4].n3 WWL[4].n2 3.576
R17445 WWL[4].n5 WWL[4].n4 3.576
R17446 WWL[4].n7 WWL[4].n6 3.576
R17447 WWL[4].n9 WWL[4].n8 3.576
R17448 WWL[4].n11 WWL[4].n10 3.576
R17449 WWL[4].n13 WWL[4].n12 3.576
R17450 WWL[4].n15 WWL[4].n14 3.576
R17451 WWL[4].n17 WWL[4].n16 3.576
R17452 WWL[4].n19 WWL[4].n18 3.576
R17453 WWL[4].n21 WWL[4].n20 3.576
R17454 WWL[4].n23 WWL[4].n22 3.576
R17455 WWL[4].n25 WWL[4].n24 3.576
R17456 WWL[4].n27 WWL[4].n26 3.576
R17457 WWL[4].n29 WWL[4].n28 3.576
R17458 WWL[4].n2 WWL[4].n1 1.317
R17459 WWL[4].n4 WWL[4].n3 1.317
R17460 WWL[4].n6 WWL[4].n5 1.317
R17461 WWL[4].n8 WWL[4].n7 1.317
R17462 WWL[4].n10 WWL[4].n9 1.317
R17463 WWL[4].n12 WWL[4].n11 1.317
R17464 WWL[4].n14 WWL[4].n13 1.317
R17465 WWL[4].n16 WWL[4].n15 1.317
R17466 WWL[4].n18 WWL[4].n17 1.317
R17467 WWL[4].n20 WWL[4].n19 1.317
R17468 WWL[4].n22 WWL[4].n21 1.317
R17469 WWL[4].n24 WWL[4].n23 1.317
R17470 WWL[4].n26 WWL[4].n25 1.317
R17471 WWL[4].n28 WWL[4].n27 1.317
R17472 WWL[4].n30 WWL[4].n29 1.317
R17473 a_5342_1939.t0 a_5342_1939.t1 242.857
R17474 a_1440_n271.t0 a_1440_n271.t1 242.857
R17475 a_n2345_n5338.n0 a_n2345_n5338.t0 63.08
R17476 a_n2345_n5338.t1 a_n2345_n5338.n0 41.303
R17477 a_n2345_n5338.n0 a_n2345_n5338.t2 2.251
R17478 a_1427_4671.n0 a_1427_4671.t2 362.857
R17479 a_1427_4671.t5 a_1427_4671.t3 337.399
R17480 a_1427_4671.t3 a_1427_4671.t4 298.839
R17481 a_1427_4671.n0 a_1427_4671.t5 280.405
R17482 a_1427_4671.n1 a_1427_4671.t0 200
R17483 a_1427_4671.n1 a_1427_4671.n0 172.311
R17484 a_1427_4671.n2 a_1427_4671.n1 24
R17485 a_1427_4671.n1 a_1427_4671.t1 21.212
R17486 a_1522_4686.n0 a_1522_4686.t2 358.166
R17487 a_1522_4686.t4 a_1522_4686.t3 337.399
R17488 a_1522_4686.t3 a_1522_4686.t5 285.986
R17489 a_1522_4686.n0 a_1522_4686.t4 282.573
R17490 a_1522_4686.n1 a_1522_4686.t0 202.857
R17491 a_1522_4686.n1 a_1522_4686.n0 173.817
R17492 a_1522_4686.n1 a_1522_4686.t1 20.826
R17493 a_1522_4686.n2 a_1522_4686.n1 20.689
R17494 a_1427_678.n0 a_1427_678.t2 362.857
R17495 a_1427_678.t4 a_1427_678.t3 337.399
R17496 a_1427_678.t3 a_1427_678.t5 298.839
R17497 a_1427_678.n0 a_1427_678.t4 280.405
R17498 a_1427_678.n1 a_1427_678.t0 200
R17499 a_1427_678.n1 a_1427_678.n0 172.311
R17500 a_1427_678.n2 a_1427_678.n1 24
R17501 a_1427_678.n1 a_1427_678.t1 21.212
R17502 a_1522_693.n0 a_1522_693.t2 358.166
R17503 a_1522_693.t5 a_1522_693.t4 337.399
R17504 a_1522_693.t4 a_1522_693.t3 285.986
R17505 a_1522_693.n0 a_1522_693.t5 282.573
R17506 a_1522_693.n1 a_1522_693.t0 202.857
R17507 a_1522_693.n1 a_1522_693.n0 173.817
R17508 a_1522_693.n1 a_1522_693.t1 20.826
R17509 a_1522_693.n2 a_1522_693.n1 20.689
R17510 a_4302_n45.n0 a_4302_n45.t1 362.857
R17511 a_4302_n45.t5 a_4302_n45.t4 337.399
R17512 a_4302_n45.t4 a_4302_n45.t3 298.839
R17513 a_4302_n45.n0 a_4302_n45.t5 280.405
R17514 a_4302_n45.n1 a_4302_n45.t2 200
R17515 a_4302_n45.n1 a_4302_n45.n0 172.311
R17516 a_4302_n45.n2 a_4302_n45.n1 24
R17517 a_4302_n45.n1 a_4302_n45.t0 21.212
R17518 a_4315_n30.t0 a_4315_n30.t1 242.857
R17519 a_8997_1939.n0 a_8997_1939.t0 358.166
R17520 a_8997_1939.t5 a_8997_1939.t3 337.399
R17521 a_8997_1939.t3 a_8997_1939.t4 285.986
R17522 a_8997_1939.n0 a_8997_1939.t5 282.573
R17523 a_8997_1939.n1 a_8997_1939.t2 202.857
R17524 a_8997_1939.n1 a_8997_1939.n0 173.817
R17525 a_8997_1939.n1 a_8997_1939.t1 20.826
R17526 a_8997_1939.n2 a_8997_1939.n1 20.689
R17527 a_8902_1924.n0 a_8902_1924.t1 362.857
R17528 a_8902_1924.t5 a_8902_1924.t4 337.399
R17529 a_8902_1924.t4 a_8902_1924.t3 298.839
R17530 a_8902_1924.n0 a_8902_1924.t5 280.405
R17531 a_8902_1924.n1 a_8902_1924.t2 200
R17532 a_8902_1924.n1 a_8902_1924.n0 172.311
R17533 a_8902_1924.n2 a_8902_1924.n1 24
R17534 a_8902_1924.n1 a_8902_1924.t0 21.212
R17535 ADC7_OUT[2].n0 ADC7_OUT[2].t4 1354.27
R17536 ADC7_OUT[2].n0 ADC7_OUT[2].t3 821.954
R17537 ADC7_OUT[2].n3 ADC7_OUT[2].t0 344.879
R17538 ADC7_OUT[2].n2 ADC7_OUT[2].t1 266.575
R17539 ADC7_OUT[2].n1 ADC7_OUT[2].n0 149.035
R17540 ADC7_OUT[2].n1 ADC7_OUT[2].t2 46.723
R17541 ADC7_OUT[2].n3 ADC7_OUT[2].n2 39.152
R17542 ADC7_OUT[2] ADC7_OUT[2].n3 38.137
R17543 ADC7_OUT[2].n2 ADC7_OUT[2].n1 17.317
R17544 a_4675_n7216.n0 a_4675_n7216.t4 1464.36
R17545 a_4675_n7216.n0 a_4675_n7216.t3 713.588
R17546 a_4675_n7216.n1 a_4675_n7216.t0 374.998
R17547 a_4675_n7216.n1 a_4675_n7216.t1 273.351
R17548 a_4675_n7216.n2 a_4675_n7216.n0 143.764
R17549 a_4675_n7216.t2 a_4675_n7216.n2 78.209
R17550 a_4675_n7216.n2 a_4675_n7216.n1 4.517
R17551 a_2853_n1770.n0 a_2853_n1770.t1 160.619
R17552 a_2853_n1770.t0 a_2853_n1770.n0 151.153
R17553 a_2660_n1770.n0 a_2660_n1770.t1 325.682
R17554 a_2660_n1770.n0 a_2660_n1770.t2 322.294
R17555 a_2660_n1770.t0 a_2660_n1770.n0 73.623
R17556 a_4972_2662.n0 a_4972_2662.t0 358.166
R17557 a_4972_2662.t3 a_4972_2662.t5 337.399
R17558 a_4972_2662.t5 a_4972_2662.t4 285.986
R17559 a_4972_2662.n0 a_4972_2662.t3 282.573
R17560 a_4972_2662.n1 a_4972_2662.t2 202.857
R17561 a_4972_2662.n1 a_4972_2662.n0 173.817
R17562 a_4972_2662.n1 a_4972_2662.t1 20.826
R17563 a_4972_2662.n2 a_4972_2662.n1 20.689
R17564 a_4877_2647.n0 a_4877_2647.t1 362.857
R17565 a_4877_2647.t4 a_4877_2647.t3 337.399
R17566 a_4877_2647.t3 a_4877_2647.t5 298.839
R17567 a_4877_2647.n0 a_4877_2647.t4 280.405
R17568 a_4877_2647.n1 a_4877_2647.t2 200
R17569 a_4877_2647.n1 a_4877_2647.n0 172.311
R17570 a_4877_2647.n2 a_4877_2647.n1 24
R17571 a_4877_2647.n1 a_4877_2647.t0 21.212
R17572 WWL[3].n0 WWL[3].t1 262.032
R17573 WWL[3].n29 WWL[3].t4 260.715
R17574 WWL[3].n27 WWL[3].t7 260.715
R17575 WWL[3].n25 WWL[3].t20 260.715
R17576 WWL[3].n23 WWL[3].t15 260.715
R17577 WWL[3].n21 WWL[3].t25 260.715
R17578 WWL[3].n19 WWL[3].t11 260.715
R17579 WWL[3].n17 WWL[3].t3 260.715
R17580 WWL[3].n15 WWL[3].t18 260.715
R17581 WWL[3].n13 WWL[3].t8 260.715
R17582 WWL[3].n11 WWL[3].t16 260.715
R17583 WWL[3].n9 WWL[3].t5 260.715
R17584 WWL[3].n7 WWL[3].t19 260.715
R17585 WWL[3].n5 WWL[3].t13 260.715
R17586 WWL[3].n3 WWL[3].t28 260.715
R17587 WWL[3].n1 WWL[3].t9 260.715
R17588 WWL[3].n30 WWL[3].t21 259.254
R17589 WWL[3].n28 WWL[3].t27 259.254
R17590 WWL[3].n26 WWL[3].t6 259.254
R17591 WWL[3].n24 WWL[3].t22 259.254
R17592 WWL[3].n22 WWL[3].t14 259.254
R17593 WWL[3].n20 WWL[3].t29 259.254
R17594 WWL[3].n18 WWL[3].t10 259.254
R17595 WWL[3].n16 WWL[3].t24 259.254
R17596 WWL[3].n14 WWL[3].t17 259.254
R17597 WWL[3].n12 WWL[3].t0 259.254
R17598 WWL[3].n10 WWL[3].t23 259.254
R17599 WWL[3].n8 WWL[3].t30 259.254
R17600 WWL[3].n6 WWL[3].t31 259.254
R17601 WWL[3].n4 WWL[3].t2 259.254
R17602 WWL[3].n2 WWL[3].t26 259.254
R17603 WWL[3].n0 WWL[3].t12 259.254
R17604 WWL[3] WWL[3].n30 44.647
R17605 WWL[3].n1 WWL[3].n0 3.576
R17606 WWL[3].n3 WWL[3].n2 3.576
R17607 WWL[3].n5 WWL[3].n4 3.576
R17608 WWL[3].n7 WWL[3].n6 3.576
R17609 WWL[3].n9 WWL[3].n8 3.576
R17610 WWL[3].n11 WWL[3].n10 3.576
R17611 WWL[3].n13 WWL[3].n12 3.576
R17612 WWL[3].n15 WWL[3].n14 3.576
R17613 WWL[3].n17 WWL[3].n16 3.576
R17614 WWL[3].n19 WWL[3].n18 3.576
R17615 WWL[3].n21 WWL[3].n20 3.576
R17616 WWL[3].n23 WWL[3].n22 3.576
R17617 WWL[3].n25 WWL[3].n24 3.576
R17618 WWL[3].n27 WWL[3].n26 3.576
R17619 WWL[3].n29 WWL[3].n28 3.576
R17620 WWL[3].n2 WWL[3].n1 1.317
R17621 WWL[3].n4 WWL[3].n3 1.317
R17622 WWL[3].n6 WWL[3].n5 1.317
R17623 WWL[3].n8 WWL[3].n7 1.317
R17624 WWL[3].n10 WWL[3].n9 1.317
R17625 WWL[3].n12 WWL[3].n11 1.317
R17626 WWL[3].n14 WWL[3].n13 1.317
R17627 WWL[3].n16 WWL[3].n15 1.317
R17628 WWL[3].n18 WWL[3].n17 1.317
R17629 WWL[3].n20 WWL[3].n19 1.317
R17630 WWL[3].n22 WWL[3].n21 1.317
R17631 WWL[3].n24 WWL[3].n23 1.317
R17632 WWL[3].n26 WWL[3].n25 1.317
R17633 WWL[3].n28 WWL[3].n27 1.317
R17634 WWL[3].n30 WWL[3].n29 1.317
R17635 a_5547_2943.n0 a_5547_2943.t1 358.166
R17636 a_5547_2943.t4 a_5547_2943.t5 337.399
R17637 a_5547_2943.t5 a_5547_2943.t3 285.986
R17638 a_5547_2943.n0 a_5547_2943.t4 282.573
R17639 a_5547_2943.n1 a_5547_2943.t2 202.857
R17640 a_5547_2943.n1 a_5547_2943.n0 173.817
R17641 a_5547_2943.n1 a_5547_2943.t0 20.826
R17642 a_5547_2943.n2 a_5547_2943.n1 20.689
R17643 RWL[9].n0 RWL[9].t12 154.243
R17644 RWL[9].n14 RWL[9].t2 149.249
R17645 RWL[9].n13 RWL[9].t7 149.249
R17646 RWL[9].n12 RWL[9].t14 149.249
R17647 RWL[9].n11 RWL[9].t3 149.249
R17648 RWL[9].n10 RWL[9].t0 149.249
R17649 RWL[9].n9 RWL[9].t8 149.249
R17650 RWL[9].n8 RWL[9].t15 149.249
R17651 RWL[9].n7 RWL[9].t5 149.249
R17652 RWL[9].n6 RWL[9].t1 149.249
R17653 RWL[9].n5 RWL[9].t11 149.249
R17654 RWL[9].n4 RWL[9].t4 149.249
R17655 RWL[9].n3 RWL[9].t9 149.249
R17656 RWL[9].n2 RWL[9].t10 149.249
R17657 RWL[9].n1 RWL[9].t13 149.249
R17658 RWL[9].n0 RWL[9].t6 149.249
R17659 RWL[9] RWL[9].n14 42.872
R17660 RWL[9].n1 RWL[9].n0 4.994
R17661 RWL[9].n2 RWL[9].n1 4.994
R17662 RWL[9].n3 RWL[9].n2 4.994
R17663 RWL[9].n4 RWL[9].n3 4.994
R17664 RWL[9].n5 RWL[9].n4 4.994
R17665 RWL[9].n6 RWL[9].n5 4.994
R17666 RWL[9].n7 RWL[9].n6 4.994
R17667 RWL[9].n8 RWL[9].n7 4.994
R17668 RWL[9].n9 RWL[9].n8 4.994
R17669 RWL[9].n10 RWL[9].n9 4.994
R17670 RWL[9].n11 RWL[9].n10 4.994
R17671 RWL[9].n12 RWL[9].n11 4.994
R17672 RWL[9].n13 RWL[9].n12 4.994
R17673 RWL[9].n14 RWL[9].n13 4.994
R17674 a_2590_1457.t0 a_2590_1457.t1 242.857
R17675 a_4877_960.n0 a_4877_960.t1 362.857
R17676 a_4877_960.t4 a_4877_960.t3 337.399
R17677 a_4877_960.t3 a_4877_960.t5 298.839
R17678 a_4877_960.n0 a_4877_960.t4 280.405
R17679 a_4877_960.n1 a_4877_960.t0 200
R17680 a_4877_960.n1 a_4877_960.n0 172.311
R17681 a_4877_960.n2 a_4877_960.n1 24
R17682 a_4877_960.n1 a_4877_960.t2 21.212
R17683 a_4877_n527.n0 a_4877_n527.t0 362.857
R17684 a_4877_n527.t4 a_4877_n527.t3 337.399
R17685 a_4877_n527.t3 a_4877_n527.t5 298.839
R17686 a_4877_n527.n0 a_4877_n527.t4 280.405
R17687 a_4877_n527.n1 a_4877_n527.t2 200
R17688 a_4877_n527.n1 a_4877_n527.n0 172.311
R17689 a_4877_n527.n2 a_4877_n527.n1 24
R17690 a_4877_n527.n1 a_4877_n527.t1 21.212
R17691 RWL[1].n0 RWL[1].t14 154.243
R17692 RWL[1].n14 RWL[1].t4 149.249
R17693 RWL[1].n13 RWL[1].t9 149.249
R17694 RWL[1].n12 RWL[1].t0 149.249
R17695 RWL[1].n11 RWL[1].t5 149.249
R17696 RWL[1].n10 RWL[1].t2 149.249
R17697 RWL[1].n9 RWL[1].t10 149.249
R17698 RWL[1].n8 RWL[1].t1 149.249
R17699 RWL[1].n7 RWL[1].t7 149.249
R17700 RWL[1].n6 RWL[1].t3 149.249
R17701 RWL[1].n5 RWL[1].t13 149.249
R17702 RWL[1].n4 RWL[1].t6 149.249
R17703 RWL[1].n3 RWL[1].t11 149.249
R17704 RWL[1].n2 RWL[1].t12 149.249
R17705 RWL[1].n1 RWL[1].t15 149.249
R17706 RWL[1].n0 RWL[1].t8 149.249
R17707 RWL[1] RWL[1].n14 42.872
R17708 RWL[1].n1 RWL[1].n0 4.994
R17709 RWL[1].n2 RWL[1].n1 4.994
R17710 RWL[1].n3 RWL[1].n2 4.994
R17711 RWL[1].n4 RWL[1].n3 4.994
R17712 RWL[1].n5 RWL[1].n4 4.994
R17713 RWL[1].n6 RWL[1].n5 4.994
R17714 RWL[1].n7 RWL[1].n6 4.994
R17715 RWL[1].n8 RWL[1].n7 4.994
R17716 RWL[1].n9 RWL[1].n8 4.994
R17717 RWL[1].n10 RWL[1].n9 4.994
R17718 RWL[1].n11 RWL[1].n10 4.994
R17719 RWL[1].n12 RWL[1].n11 4.994
R17720 RWL[1].n13 RWL[1].n12 4.994
R17721 RWL[1].n14 RWL[1].n13 4.994
R17722 a_1440_3425.t0 a_1440_3425.t1 242.857
R17723 a_1050_n2132.n0 a_1050_n2132.t2 489.336
R17724 a_1050_n2132.n0 a_1050_n2132.t1 243.258
R17725 a_1050_n2132.t0 a_1050_n2132.n0 214.415
R17726 a_8997_2662.n0 a_8997_2662.t1 358.166
R17727 a_8997_2662.t4 a_8997_2662.t5 337.399
R17728 a_8997_2662.t5 a_8997_2662.t3 285.986
R17729 a_8997_2662.n0 a_8997_2662.t4 282.573
R17730 a_8997_2662.n1 a_8997_2662.t2 202.857
R17731 a_8997_2662.n1 a_8997_2662.n0 173.817
R17732 a_8997_2662.n1 a_8997_2662.t0 20.826
R17733 a_8997_2662.n2 a_8997_2662.n1 20.689
R17734 a_9367_2662.t0 a_9367_2662.t1 242.857
R17735 a_5342_1698.t0 a_5342_1698.t1 242.857
R17736 a_1892_693.t0 a_1892_693.t1 242.857
R17737 ADC1_OUT[1].n0 ADC1_OUT[1].t4 1355.37
R17738 ADC1_OUT[1].n0 ADC1_OUT[1].t3 820.859
R17739 ADC1_OUT[1].n3 ADC1_OUT[1].t0 336.667
R17740 ADC1_OUT[1].n2 ADC1_OUT[1].t2 266.644
R17741 ADC1_OUT[1].n1 ADC1_OUT[1].n0 149.035
R17742 ADC1_OUT[1].n3 ADC1_OUT[1].n2 47.435
R17743 ADC1_OUT[1].n1 ADC1_OUT[1].t1 45.968
R17744 ADC1_OUT[1] ADC1_OUT[1].n3 45.936
R17745 ADC1_OUT[1].n2 ADC1_OUT[1].n1 17.317
R17746 a_n2642_n5293.n0 a_n2642_n5293.t0 65.063
R17747 a_n2642_n5293.n0 a_n2642_n5293.t2 42.011
R17748 a_n2642_n5293.t1 a_n2642_n5293.n0 2.113
R17749 RWLB[13].n0 RWLB[13].t1 154.228
R17750 RWLB[13].n14 RWLB[13].t6 149.249
R17751 RWLB[13].n13 RWLB[13].t5 149.249
R17752 RWLB[13].n12 RWLB[13].t13 149.249
R17753 RWLB[13].n11 RWLB[13].t9 149.249
R17754 RWLB[13].n10 RWLB[13].t0 149.249
R17755 RWLB[13].n9 RWLB[13].t15 149.249
R17756 RWLB[13].n8 RWLB[13].t3 149.249
R17757 RWLB[13].n7 RWLB[13].t2 149.249
R17758 RWLB[13].n6 RWLB[13].t11 149.249
R17759 RWLB[13].n5 RWLB[13].t10 149.249
R17760 RWLB[13].n4 RWLB[13].t12 149.249
R17761 RWLB[13].n3 RWLB[13].t7 149.249
R17762 RWLB[13].n2 RWLB[13].t4 149.249
R17763 RWLB[13].n1 RWLB[13].t14 149.249
R17764 RWLB[13].n0 RWLB[13].t8 149.249
R17765 RWLB[13] RWLB[13].n14 47.816
R17766 RWLB[13].n1 RWLB[13].n0 4.979
R17767 RWLB[13].n2 RWLB[13].n1 4.979
R17768 RWLB[13].n3 RWLB[13].n2 4.979
R17769 RWLB[13].n4 RWLB[13].n3 4.979
R17770 RWLB[13].n5 RWLB[13].n4 4.979
R17771 RWLB[13].n6 RWLB[13].n5 4.979
R17772 RWLB[13].n7 RWLB[13].n6 4.979
R17773 RWLB[13].n8 RWLB[13].n7 4.979
R17774 RWLB[13].n9 RWLB[13].n8 4.979
R17775 RWLB[13].n10 RWLB[13].n9 4.979
R17776 RWLB[13].n11 RWLB[13].n10 4.979
R17777 RWLB[13].n12 RWLB[13].n11 4.979
R17778 RWLB[13].n13 RWLB[13].n12 4.979
R17779 RWLB[13].n14 RWLB[13].n13 4.979
R17780 a_3042_452.t0 a_3042_452.t1 242.857
R17781 a_7752_4671.n0 a_7752_4671.t2 362.857
R17782 a_7752_4671.t4 a_7752_4671.t5 337.399
R17783 a_7752_4671.t5 a_7752_4671.t3 298.839
R17784 a_7752_4671.n0 a_7752_4671.t4 280.405
R17785 a_7752_4671.n1 a_7752_4671.t0 200
R17786 a_7752_4671.n1 a_7752_4671.n0 172.311
R17787 a_7752_4671.n2 a_7752_4671.n1 24
R17788 a_7752_4671.n1 a_7752_4671.t1 21.212
R17789 a_7765_4686.t0 a_7765_4686.t1 242.857
R17790 WWL[6].n0 WWL[6].t9 262.032
R17791 WWL[6].n29 WWL[6].t12 260.715
R17792 WWL[6].n27 WWL[6].t15 260.715
R17793 WWL[6].n25 WWL[6].t29 260.715
R17794 WWL[6].n23 WWL[6].t23 260.715
R17795 WWL[6].n21 WWL[6].t3 260.715
R17796 WWL[6].n19 WWL[6].t20 260.715
R17797 WWL[6].n17 WWL[6].t11 260.715
R17798 WWL[6].n15 WWL[6].t26 260.715
R17799 WWL[6].n13 WWL[6].t16 260.715
R17800 WWL[6].n11 WWL[6].t24 260.715
R17801 WWL[6].n9 WWL[6].t13 260.715
R17802 WWL[6].n7 WWL[6].t27 260.715
R17803 WWL[6].n5 WWL[6].t21 260.715
R17804 WWL[6].n3 WWL[6].t4 260.715
R17805 WWL[6].n1 WWL[6].t17 260.715
R17806 WWL[6].n30 WWL[6].t28 259.254
R17807 WWL[6].n28 WWL[6].t2 259.254
R17808 WWL[6].n26 WWL[6].t14 259.254
R17809 WWL[6].n24 WWL[6].t30 259.254
R17810 WWL[6].n22 WWL[6].t22 259.254
R17811 WWL[6].n20 WWL[6].t5 259.254
R17812 WWL[6].n18 WWL[6].t18 259.254
R17813 WWL[6].n16 WWL[6].t0 259.254
R17814 WWL[6].n14 WWL[6].t25 259.254
R17815 WWL[6].n12 WWL[6].t8 259.254
R17816 WWL[6].n10 WWL[6].t31 259.254
R17817 WWL[6].n8 WWL[6].t6 259.254
R17818 WWL[6].n6 WWL[6].t7 259.254
R17819 WWL[6].n4 WWL[6].t10 259.254
R17820 WWL[6].n2 WWL[6].t1 259.254
R17821 WWL[6].n0 WWL[6].t19 259.254
R17822 WWL[6] WWL[6].n30 44.647
R17823 WWL[6].n1 WWL[6].n0 3.576
R17824 WWL[6].n3 WWL[6].n2 3.576
R17825 WWL[6].n5 WWL[6].n4 3.576
R17826 WWL[6].n7 WWL[6].n6 3.576
R17827 WWL[6].n9 WWL[6].n8 3.576
R17828 WWL[6].n11 WWL[6].n10 3.576
R17829 WWL[6].n13 WWL[6].n12 3.576
R17830 WWL[6].n15 WWL[6].n14 3.576
R17831 WWL[6].n17 WWL[6].n16 3.576
R17832 WWL[6].n19 WWL[6].n18 3.576
R17833 WWL[6].n21 WWL[6].n20 3.576
R17834 WWL[6].n23 WWL[6].n22 3.576
R17835 WWL[6].n25 WWL[6].n24 3.576
R17836 WWL[6].n27 WWL[6].n26 3.576
R17837 WWL[6].n29 WWL[6].n28 3.576
R17838 WWL[6].n2 WWL[6].n1 1.317
R17839 WWL[6].n4 WWL[6].n3 1.317
R17840 WWL[6].n6 WWL[6].n5 1.317
R17841 WWL[6].n8 WWL[6].n7 1.317
R17842 WWL[6].n10 WWL[6].n9 1.317
R17843 WWL[6].n12 WWL[6].n11 1.317
R17844 WWL[6].n14 WWL[6].n13 1.317
R17845 WWL[6].n16 WWL[6].n15 1.317
R17846 WWL[6].n18 WWL[6].n17 1.317
R17847 WWL[6].n20 WWL[6].n19 1.317
R17848 WWL[6].n22 WWL[6].n21 1.317
R17849 WWL[6].n24 WWL[6].n23 1.317
R17850 WWL[6].n26 WWL[6].n25 1.317
R17851 WWL[6].n28 WWL[6].n27 1.317
R17852 WWL[6].n30 WWL[6].n29 1.317
R17853 a_6615_1698.t0 a_6615_1698.t1 242.857
R17854 a_10856_n4114.t1 a_10856_n4114.t0 336.812
R17855 a_2577_437.n0 a_2577_437.t0 362.857
R17856 a_2577_437.t3 a_2577_437.t5 337.399
R17857 a_2577_437.t5 a_2577_437.t4 298.839
R17858 a_2577_437.n0 a_2577_437.t3 280.405
R17859 a_2577_437.n1 a_2577_437.t2 200
R17860 a_2577_437.n1 a_2577_437.n0 172.311
R17861 a_2577_437.n2 a_2577_437.n1 24
R17862 a_2577_437.n1 a_2577_437.t1 21.212
R17863 a_2672_452.n0 a_2672_452.t1 358.166
R17864 a_2672_452.t4 a_2672_452.t3 337.399
R17865 a_2672_452.t3 a_2672_452.t5 285.986
R17866 a_2672_452.n0 a_2672_452.t4 282.573
R17867 a_2672_452.n1 a_2672_452.t2 202.857
R17868 a_2672_452.n1 a_2672_452.n0 173.817
R17869 a_2672_452.n1 a_2672_452.t0 20.826
R17870 a_2672_452.n2 a_2672_452.n1 20.689
R17871 Iref2.n0 Iref2.t7 463.323
R17872 Iref2.n14 Iref2.t6 454.171
R17873 Iref2.n13 Iref2.t15 454.171
R17874 Iref2.n12 Iref2.t8 454.171
R17875 Iref2.n11 Iref2.t14 454.171
R17876 Iref2.n10 Iref2.t13 454.171
R17877 Iref2.n9 Iref2.t1 454.171
R17878 Iref2.n8 Iref2.t4 454.171
R17879 Iref2.n7 Iref2.t11 454.171
R17880 Iref2.n6 Iref2.t3 454.171
R17881 Iref2.n5 Iref2.t10 454.171
R17882 Iref2.n4 Iref2.t2 454.171
R17883 Iref2.n3 Iref2.t9 454.171
R17884 Iref2.n2 Iref2.t12 454.171
R17885 Iref2.n1 Iref2.t5 454.171
R17886 Iref2.n0 Iref2.t0 454.171
R17887 Iref2 Iref2.n14 20.357
R17888 Iref2.n12 Iref2.n11 8.671
R17889 Iref2.n13 Iref2.n12 8.671
R17890 Iref2.n10 Iref2.n9 8.649
R17891 Iref2.n11 Iref2.n10 8.649
R17892 Iref2.n1 Iref2.n0 8.634
R17893 Iref2.n4 Iref2.n3 8.634
R17894 Iref2.n5 Iref2.n4 8.634
R17895 Iref2.n6 Iref2.n5 8.634
R17896 Iref2.n7 Iref2.n6 8.634
R17897 Iref2.n8 Iref2.n7 8.634
R17898 Iref2.n9 Iref2.n8 8.634
R17899 Iref2.n2 Iref2.n1 8.627
R17900 Iref2.n3 Iref2.n2 8.627
R17901 Iref2.n14 Iref2.n13 6.568
R17902 a_n2148_n6847.t1 a_n2148_n6847.t0 336.812
R17903 a_n2207_n7203.t0 a_n2207_n7203.t1 68.741
R17904 a_5857_n7216.n0 a_5857_n7216.t3 1464.36
R17905 a_5857_n7216.n0 a_5857_n7216.t4 713.588
R17906 a_5857_n7216.n1 a_5857_n7216.t0 374.998
R17907 a_5857_n7216.n1 a_5857_n7216.t2 273.351
R17908 a_5857_n7216.n2 a_5857_n7216.n0 143.764
R17909 a_5857_n7216.t1 a_5857_n7216.n2 78.209
R17910 a_5857_n7216.n2 a_5857_n7216.n1 4.517
R17911 a_5630_n6503.n0 a_5630_n6503.t0 65.064
R17912 a_5630_n6503.n0 a_5630_n6503.t2 42.011
R17913 a_5630_n6503.t1 a_5630_n6503.n0 2.113
R17914 a_6812_n3770.n0 a_6812_n3770.t0 65.064
R17915 a_6812_n3770.t1 a_6812_n3770.n0 42.011
R17916 a_6812_n3770.n0 a_6812_n3770.t2 2.113
R17917 a_3165_1216.t0 a_3165_1216.t1 242.857
R17918 a_6027_1201.n0 a_6027_1201.t1 362.857
R17919 a_6027_1201.t5 a_6027_1201.t3 337.399
R17920 a_6027_1201.t3 a_6027_1201.t4 298.839
R17921 a_6027_1201.n0 a_6027_1201.t5 280.405
R17922 a_6027_1201.n1 a_6027_1201.t0 200
R17923 a_6027_1201.n1 a_6027_1201.n0 172.311
R17924 a_6027_1201.n2 a_6027_1201.n1 24
R17925 a_6027_1201.n1 a_6027_1201.t2 21.212
R17926 a_6122_1216.n0 a_6122_1216.t2 358.166
R17927 a_6122_1216.t4 a_6122_1216.t3 337.399
R17928 a_6122_1216.t3 a_6122_1216.t5 285.986
R17929 a_6122_1216.n0 a_6122_1216.t4 282.573
R17930 a_6122_1216.n1 a_6122_1216.t0 202.857
R17931 a_6122_1216.n1 a_6122_1216.n0 173.817
R17932 a_6122_1216.n1 a_6122_1216.t1 20.826
R17933 a_6122_1216.n2 a_6122_1216.n1 20.689
R17934 a_5728_n1770.n0 a_5728_n1770.t1 160.619
R17935 a_5728_n1770.t0 a_5728_n1770.n0 151.153
R17936 a_5535_n1770.n0 a_5535_n1770.t2 322.294
R17937 a_5535_n1770.n1 a_5535_n1770.n0 229.466
R17938 a_5535_n1770.t0 a_5535_n1770.n1 151.15
R17939 a_5535_n1770.n0 a_5535_n1770.t1 73.623
R17940 a_6615_n812.t0 a_6615_n812.t1 242.857
R17941 ADC8_OUT[0].n0 ADC8_OUT[0].t4 1354.27
R17942 ADC8_OUT[0].n0 ADC8_OUT[0].t3 821.954
R17943 ADC8_OUT[0].n3 ADC8_OUT[0].t0 341.115
R17944 ADC8_OUT[0].n2 ADC8_OUT[0].t2 266.575
R17945 ADC8_OUT[0].n1 ADC8_OUT[0].n0 149.035
R17946 ADC8_OUT[0] ADC8_OUT[0].n3 61.811
R17947 ADC8_OUT[0].n1 ADC8_OUT[0].t1 46.723
R17948 ADC8_OUT[0].n3 ADC8_OUT[0].n2 42.917
R17949 ADC8_OUT[0].n2 ADC8_OUT[0].n1 17.317
R17950 a_5857_n4483.n0 a_5857_n4483.t3 1464.36
R17951 a_5857_n4483.n0 a_5857_n4483.t4 713.588
R17952 a_5857_n4483.n1 a_5857_n4483.t0 374.998
R17953 a_5857_n4483.n1 a_5857_n4483.t2 273.351
R17954 a_5857_n4483.n2 a_5857_n4483.n0 143.764
R17955 a_5857_n4483.t1 a_5857_n4483.n2 78.209
R17956 a_5857_n4483.n2 a_5857_n4483.n1 4.517
R17957 a_n3565_n7216.n0 a_n3565_n7216.t4 1464.36
R17958 a_n3565_n7216.n0 a_n3565_n7216.t3 713.588
R17959 a_n3565_n7216.n1 a_n3565_n7216.t0 374.998
R17960 a_n3565_n7216.n1 a_n3565_n7216.t1 273.351
R17961 a_n3565_n7216.n2 a_n3565_n7216.n0 143.764
R17962 a_n3565_n7216.t2 a_n3565_n7216.n2 78.209
R17963 a_n3565_n7216.n2 a_n3565_n7216.n1 4.517
R17964 a_7994_n6503.n0 a_7994_n6503.t0 65.064
R17965 a_7994_n6503.n0 a_7994_n6503.t2 42.011
R17966 a_7994_n6503.t1 a_7994_n6503.n0 2.113
R17967 a_1427_2165.n0 a_1427_2165.t1 362.857
R17968 a_1427_2165.t3 a_1427_2165.t4 337.399
R17969 a_1427_2165.t4 a_1427_2165.t5 298.839
R17970 a_1427_2165.n0 a_1427_2165.t3 280.405
R17971 a_1427_2165.n1 a_1427_2165.t0 200
R17972 a_1427_2165.n1 a_1427_2165.n0 172.311
R17973 a_1427_2165.n2 a_1427_2165.n1 24
R17974 a_1427_2165.n1 a_1427_2165.t2 21.212
R17975 a_1522_2180.n0 a_1522_2180.t2 358.166
R17976 a_1522_2180.t5 a_1522_2180.t4 337.399
R17977 a_1522_2180.t4 a_1522_2180.t3 285.986
R17978 a_1522_2180.n0 a_1522_2180.t5 282.573
R17979 a_1522_2180.n1 a_1522_2180.t0 202.857
R17980 a_1522_2180.n1 a_1522_2180.n0 173.817
R17981 a_1522_2180.n1 a_1522_2180.t1 20.826
R17982 a_1522_2180.n2 a_1522_2180.n1 20.689
R17983 ADC12_OUT[2].n0 ADC12_OUT[2].t4 1354.27
R17984 ADC12_OUT[2].n0 ADC12_OUT[2].t3 821.954
R17985 ADC12_OUT[2].n3 ADC12_OUT[2].t0 333.585
R17986 ADC12_OUT[2].n2 ADC12_OUT[2].t2 266.575
R17987 ADC12_OUT[2].n1 ADC12_OUT[2].n0 149.035
R17988 ADC12_OUT[2].n3 ADC12_OUT[2].n2 50.447
R17989 ADC12_OUT[2].n1 ADC12_OUT[2].t1 46.723
R17990 ADC12_OUT[2] ADC12_OUT[2].n3 38.164
R17991 ADC12_OUT[2].n2 ADC12_OUT[2].n1 17.317
R17992 a_3802_n2234.n2 a_3802_n2234.t1 282.97
R17993 a_3802_n2234.n1 a_3802_n2234.t3 240.683
R17994 a_3802_n2234.n0 a_3802_n2234.t4 209.208
R17995 a_3802_n2234.n0 a_3802_n2234.t2 194.167
R17996 a_3802_n2234.t0 a_3802_n2234.n2 183.404
R17997 a_3802_n2234.n1 a_3802_n2234.n0 14.805
R17998 a_3802_n2234.n2 a_3802_n2234.n1 6.415
R17999 a_3925_n2132.n0 a_3925_n2132.t2 489.336
R18000 a_3925_n2132.n0 a_3925_n2132.t1 243.258
R18001 a_3925_n2132.t0 a_3925_n2132.n0 214.415
R18002 a_8422_2421.n0 a_8422_2421.t1 358.166
R18003 a_8422_2421.t5 a_8422_2421.t4 337.399
R18004 a_8422_2421.t4 a_8422_2421.t3 285.986
R18005 a_8422_2421.n0 a_8422_2421.t5 282.573
R18006 a_8422_2421.n1 a_8422_2421.t0 202.857
R18007 a_8422_2421.n1 a_8422_2421.n0 173.817
R18008 a_8422_2421.n1 a_8422_2421.t2 20.826
R18009 a_8422_2421.n2 a_8422_2421.n1 20.689
R18010 a_8792_2421.t0 a_8792_2421.t1 242.857
R18011 a_3247_1698.n0 a_3247_1698.t0 358.166
R18012 a_3247_1698.t5 a_3247_1698.t3 337.399
R18013 a_3247_1698.t3 a_3247_1698.t4 285.986
R18014 a_3247_1698.n0 a_3247_1698.t5 282.573
R18015 a_3247_1698.n1 a_3247_1698.t2 202.857
R18016 a_3247_1698.n1 a_3247_1698.n0 173.817
R18017 a_3247_1698.n1 a_3247_1698.t1 20.826
R18018 a_3247_1698.n2 a_3247_1698.n1 20.689
R18019 a_3152_1683.n0 a_3152_1683.t1 362.857
R18020 a_3152_1683.t3 a_3152_1683.t4 337.399
R18021 a_3152_1683.t4 a_3152_1683.t5 298.839
R18022 a_3152_1683.n0 a_3152_1683.t3 280.405
R18023 a_3152_1683.n1 a_3152_1683.t2 200
R18024 a_3152_1683.n1 a_3152_1683.n0 172.311
R18025 a_3152_1683.n2 a_3152_1683.n1 24
R18026 a_3152_1683.n1 a_3152_1683.t0 21.212
R18027 ADC4_OUT[0].n0 ADC4_OUT[0].t3 1354.27
R18028 ADC4_OUT[0].n0 ADC4_OUT[0].t4 821.954
R18029 ADC4_OUT[0].n3 ADC4_OUT[0].t0 347.891
R18030 ADC4_OUT[0].n2 ADC4_OUT[0].t1 266.575
R18031 ADC4_OUT[0].n1 ADC4_OUT[0].n0 149.035
R18032 ADC4_OUT[0] ADC4_OUT[0].n3 61.508
R18033 ADC4_OUT[0].n1 ADC4_OUT[0].t2 46.723
R18034 ADC4_OUT[0].n3 ADC4_OUT[0].n2 36.141
R18035 ADC4_OUT[0].n2 ADC4_OUT[0].n1 17.317
R18036 a_3822_1939.n0 a_3822_1939.t1 358.166
R18037 a_3822_1939.t5 a_3822_1939.t4 337.399
R18038 a_3822_1939.t4 a_3822_1939.t3 285.986
R18039 a_3822_1939.n0 a_3822_1939.t5 282.573
R18040 a_3822_1939.n1 a_3822_1939.t2 202.857
R18041 a_3822_1939.n1 a_3822_1939.n0 173.817
R18042 a_3822_1939.n1 a_3822_1939.t0 20.826
R18043 a_3822_1939.n2 a_3822_1939.n1 20.689
R18044 a_3833_n953.n25 a_3833_n953.t27 561.971
R18045 a_3833_n953.n0 a_3833_n953.t5 461.908
R18046 a_3833_n953.t14 a_3833_n953.n25 108.635
R18047 a_3833_n953.n0 a_3833_n953.t6 79.512
R18048 a_3833_n953.n24 a_3833_n953.t20 65.401
R18049 a_3833_n953.n23 a_3833_n953.t1 65.401
R18050 a_3833_n953.n22 a_3833_n953.t13 65.401
R18051 a_3833_n953.n21 a_3833_n953.t15 65.401
R18052 a_3833_n953.n20 a_3833_n953.t22 65.401
R18053 a_3833_n953.n19 a_3833_n953.t18 65.401
R18054 a_3833_n953.n18 a_3833_n953.t19 65.401
R18055 a_3833_n953.n17 a_3833_n953.t10 65.401
R18056 a_3833_n953.n16 a_3833_n953.t4 65.401
R18057 a_3833_n953.n15 a_3833_n953.t8 65.401
R18058 a_3833_n953.n14 a_3833_n953.t21 65.401
R18059 a_3833_n953.n13 a_3833_n953.t23 65.401
R18060 a_3833_n953.n12 a_3833_n953.t17 65.401
R18061 a_3833_n953.n11 a_3833_n953.t11 65.401
R18062 a_3833_n953.n10 a_3833_n953.t12 65.401
R18063 a_3833_n953.n9 a_3833_n953.t24 65.401
R18064 a_3833_n953.n8 a_3833_n953.t0 65.401
R18065 a_3833_n953.n7 a_3833_n953.t3 65.401
R18066 a_3833_n953.n6 a_3833_n953.t2 65.401
R18067 a_3833_n953.n5 a_3833_n953.t26 65.401
R18068 a_3833_n953.n4 a_3833_n953.t9 65.401
R18069 a_3833_n953.n3 a_3833_n953.t16 65.401
R18070 a_3833_n953.n2 a_3833_n953.t25 65.401
R18071 a_3833_n953.n1 a_3833_n953.t7 65.401
R18072 a_3833_n953.n1 a_3833_n953.n0 5.64
R18073 a_3833_n953.n25 a_3833_n953.n24 4.438
R18074 a_3833_n953.n23 a_3833_n953.n22 2.524
R18075 a_3833_n953.n3 a_3833_n953.n2 2.498
R18076 a_3833_n953.n17 a_3833_n953.n16 2.364
R18077 a_3833_n953.n9 a_3833_n953.n8 2.355
R18078 a_3833_n953.n2 a_3833_n953.n1 1.998
R18079 a_3833_n953.n4 a_3833_n953.n3 1.998
R18080 a_3833_n953.n5 a_3833_n953.n4 1.998
R18081 a_3833_n953.n6 a_3833_n953.n5 1.998
R18082 a_3833_n953.n7 a_3833_n953.n6 1.998
R18083 a_3833_n953.n8 a_3833_n953.n7 1.998
R18084 a_3833_n953.n10 a_3833_n953.n9 1.998
R18085 a_3833_n953.n11 a_3833_n953.n10 1.998
R18086 a_3833_n953.n12 a_3833_n953.n11 1.998
R18087 a_3833_n953.n13 a_3833_n953.n12 1.998
R18088 a_3833_n953.n14 a_3833_n953.n13 1.998
R18089 a_3833_n953.n15 a_3833_n953.n14 1.998
R18090 a_3833_n953.n16 a_3833_n953.n15 1.998
R18091 a_3833_n953.n18 a_3833_n953.n17 1.998
R18092 a_3833_n953.n19 a_3833_n953.n18 1.998
R18093 a_3833_n953.n20 a_3833_n953.n19 1.998
R18094 a_3833_n953.n21 a_3833_n953.n20 1.998
R18095 a_3833_n953.n22 a_3833_n953.n21 1.998
R18096 a_3833_n953.n24 a_3833_n953.n23 1.998
R18097 a_8217_975.t0 a_8217_975.t1 242.857
R18098 a_8327_n527.n0 a_8327_n527.t1 362.857
R18099 a_8327_n527.t3 a_8327_n527.t4 337.399
R18100 a_8327_n527.t4 a_8327_n527.t5 298.839
R18101 a_8327_n527.n0 a_8327_n527.t3 280.405
R18102 a_8327_n527.n1 a_8327_n527.t2 200
R18103 a_8327_n527.n1 a_8327_n527.n0 172.311
R18104 a_8327_n527.n2 a_8327_n527.n1 24
R18105 a_8327_n527.n1 a_8327_n527.t0 21.212
R18106 a_1317_4445.t0 a_1317_4445.t1 242.857
R18107 a_6697_4148.n0 a_6697_4148.t1 358.166
R18108 a_6697_4148.t3 a_6697_4148.t4 337.399
R18109 a_6697_4148.t4 a_6697_4148.t5 285.986
R18110 a_6697_4148.n0 a_6697_4148.t3 282.573
R18111 a_6697_4148.n1 a_6697_4148.t2 202.857
R18112 a_6697_4148.n1 a_6697_4148.n0 173.817
R18113 a_6697_4148.n1 a_6697_4148.t0 20.826
R18114 a_6697_4148.n2 a_6697_4148.n1 20.689
R18115 a_3247_n812.n0 a_3247_n812.t1 358.166
R18116 a_3247_n812.t5 a_3247_n812.t3 337.399
R18117 a_3247_n812.t3 a_3247_n812.t4 285.986
R18118 a_3247_n812.n0 a_3247_n812.t5 282.573
R18119 a_3247_n812.n1 a_3247_n812.t0 202.857
R18120 a_3247_n812.n1 a_3247_n812.n0 173.817
R18121 a_3247_n812.n1 a_3247_n812.t2 20.826
R18122 a_3247_n812.n2 a_3247_n812.n1 20.689
R18123 a_3152_n827.n0 a_3152_n827.t2 362.857
R18124 a_3152_n827.t3 a_3152_n827.t4 337.399
R18125 a_3152_n827.t4 a_3152_n827.t5 298.839
R18126 a_3152_n827.n0 a_3152_n827.t3 280.405
R18127 a_3152_n827.n1 a_3152_n827.t0 200
R18128 a_3152_n827.n1 a_3152_n827.n0 172.311
R18129 a_3152_n827.n2 a_3152_n827.n1 24
R18130 a_3152_n827.n1 a_3152_n827.t1 21.212
R18131 a_9143_n4116.t0 a_9143_n4116.t1 42.707
R18132 a_9178_n3770.n0 a_9178_n3770.t0 65.064
R18133 a_9178_n3770.n0 a_9178_n3770.t2 42.011
R18134 a_9178_n3770.t1 a_9178_n3770.n0 2.113
R18135 a_1522_3907.n0 a_1522_3907.t2 358.166
R18136 a_1522_3907.t5 a_1522_3907.t4 337.399
R18137 a_1522_3907.t4 a_1522_3907.t3 285.986
R18138 a_1522_3907.n0 a_1522_3907.t5 282.573
R18139 a_1522_3907.n1 a_1522_3907.t0 202.857
R18140 a_1522_3907.n1 a_1522_3907.n0 173.817
R18141 a_1522_3907.n1 a_1522_3907.t1 20.826
R18142 a_1522_3907.n2 a_1522_3907.n1 20.689
R18143 a_1892_3907.t0 a_1892_3907.t1 242.857
R18144 a_5342_1216.t0 a_5342_1216.t1 242.857
R18145 a_2077_n2234.n2 a_2077_n2234.t0 282.97
R18146 a_2077_n2234.n1 a_2077_n2234.t3 240.683
R18147 a_2077_n2234.n0 a_2077_n2234.t4 209.208
R18148 a_2077_n2234.n0 a_2077_n2234.t2 194.167
R18149 a_2077_n2234.t1 a_2077_n2234.n2 183.404
R18150 a_2077_n2234.n1 a_2077_n2234.n0 14.805
R18151 a_2077_n2234.n2 a_2077_n2234.n1 6.415
R18152 a_2200_n2132.n0 a_2200_n2132.t2 489.336
R18153 a_2200_n2132.n0 a_2200_n2132.t1 243.258
R18154 a_2200_n2132.t0 a_2200_n2132.n0 214.415
R18155 a_2002_3651.n0 a_2002_3651.t0 362.857
R18156 a_2002_3651.t3 a_2002_3651.t5 337.399
R18157 a_2002_3651.t5 a_2002_3651.t4 298.839
R18158 a_2002_3651.n0 a_2002_3651.t3 280.405
R18159 a_2002_3651.n1 a_2002_3651.t2 200
R18160 a_2002_3651.n1 a_2002_3651.n0 172.311
R18161 a_2002_3651.n2 a_2002_3651.n1 24
R18162 a_2002_3651.n1 a_2002_3651.t1 21.212
R18163 a_7847_2662.n0 a_7847_2662.t0 358.166
R18164 a_7847_2662.t5 a_7847_2662.t3 337.399
R18165 a_7847_2662.t3 a_7847_2662.t4 285.986
R18166 a_7847_2662.n0 a_7847_2662.t5 282.573
R18167 a_7847_2662.n1 a_7847_2662.t2 202.857
R18168 a_7847_2662.n1 a_7847_2662.n0 173.817
R18169 a_7847_2662.n1 a_7847_2662.t1 20.826
R18170 a_7847_2662.n2 a_7847_2662.n1 20.689
R18171 a_4302_196.n0 a_4302_196.t2 362.857
R18172 a_4302_196.t4 a_4302_196.t3 337.399
R18173 a_4302_196.t3 a_4302_196.t5 298.839
R18174 a_4302_196.n0 a_4302_196.t4 280.405
R18175 a_4302_196.n1 a_4302_196.t1 200
R18176 a_4302_196.n1 a_4302_196.n0 172.311
R18177 a_4302_196.n2 a_4302_196.n1 24
R18178 a_4302_196.n1 a_4302_196.t0 21.212
R18179 a_7847_n30.n0 a_7847_n30.t0 358.166
R18180 a_7847_n30.t3 a_7847_n30.t5 337.399
R18181 a_7847_n30.t5 a_7847_n30.t4 285.986
R18182 a_7847_n30.n0 a_7847_n30.t3 282.573
R18183 a_7847_n30.n1 a_7847_n30.t1 202.857
R18184 a_7847_n30.n1 a_7847_n30.n0 173.817
R18185 a_7847_n30.n1 a_7847_n30.t2 20.826
R18186 a_7847_n30.n2 a_7847_n30.n1 20.689
R18187 a_7752_n45.n0 a_7752_n45.t2 362.857
R18188 a_7752_n45.t4 a_7752_n45.t3 337.399
R18189 a_7752_n45.t3 a_7752_n45.t5 298.839
R18190 a_7752_n45.n0 a_7752_n45.t4 280.405
R18191 a_7752_n45.n1 a_7752_n45.t0 200
R18192 a_7752_n45.n1 a_7752_n45.n0 172.311
R18193 a_7752_n45.n2 a_7752_n45.n1 24
R18194 a_7752_n45.n1 a_7752_n45.t1 21.212
R18195 a_5465_n512.t0 a_5465_n512.t1 242.857
R18196 a_6040_3666.t0 a_6040_3666.t1 242.857
R18197 a_7190_1698.t0 a_7190_1698.t1 242.857
R18198 a_2672_1457.n0 a_2672_1457.t2 358.166
R18199 a_2672_1457.t5 a_2672_1457.t3 337.399
R18200 a_2672_1457.t3 a_2672_1457.t4 285.986
R18201 a_2672_1457.n0 a_2672_1457.t5 282.573
R18202 a_2672_1457.n1 a_2672_1457.t0 202.857
R18203 a_2672_1457.n1 a_2672_1457.n0 173.817
R18204 a_2672_1457.n1 a_2672_1457.t1 20.826
R18205 a_2672_1457.n2 a_2672_1457.n1 20.689
R18206 a_2577_1442.n0 a_2577_1442.t2 362.857
R18207 a_2577_1442.t5 a_2577_1442.t3 337.399
R18208 a_2577_1442.t3 a_2577_1442.t4 298.839
R18209 a_2577_1442.n0 a_2577_1442.t5 280.405
R18210 a_2577_1442.n1 a_2577_1442.t0 200
R18211 a_2577_1442.n1 a_2577_1442.n0 172.311
R18212 a_2577_1442.n2 a_2577_1442.n1 24
R18213 a_2577_1442.n1 a_2577_1442.t1 21.212
R18214 a_6615_1216.t0 a_6615_1216.t1 242.857
R18215 a_n52_n4483.n0 a_n52_n4483.t3 1464.36
R18216 a_n52_n4483.n0 a_n52_n4483.t4 713.588
R18217 a_n52_n4483.n1 a_n52_n4483.t0 374.998
R18218 a_n52_n4483.n1 a_n52_n4483.t2 273.351
R18219 a_n52_n4483.n2 a_n52_n4483.n0 143.764
R18220 a_n52_n4483.t1 a_n52_n4483.n2 78.209
R18221 a_n52_n4483.n2 a_n52_n4483.n1 4.517
R18222 ADC3_OUT[0].n0 ADC3_OUT[0].t3 1354.27
R18223 ADC3_OUT[0].n0 ADC3_OUT[0].t4 821.954
R18224 ADC3_OUT[0].n3 ADC3_OUT[0].t0 344.126
R18225 ADC3_OUT[0].n2 ADC3_OUT[0].t1 266.575
R18226 ADC3_OUT[0].n1 ADC3_OUT[0].n0 149.035
R18227 ADC3_OUT[0] ADC3_OUT[0].n3 61.436
R18228 ADC3_OUT[0].n1 ADC3_OUT[0].t2 46.723
R18229 ADC3_OUT[0].n3 ADC3_OUT[0].n2 39.905
R18230 ADC3_OUT[0].n2 ADC3_OUT[0].n1 17.317
R18231 a_n279_n3770.n0 a_n279_n3770.t0 65.064
R18232 a_n279_n3770.n0 a_n279_n3770.t2 42.011
R18233 a_n279_n3770.t1 a_n279_n3770.n0 2.113
R18234 a_8422_1939.n0 a_8422_1939.t2 358.166
R18235 a_8422_1939.t3 a_8422_1939.t5 337.399
R18236 a_8422_1939.t5 a_8422_1939.t4 285.986
R18237 a_8422_1939.n0 a_8422_1939.t3 282.573
R18238 a_8422_1939.n1 a_8422_1939.t0 202.857
R18239 a_8422_1939.n1 a_8422_1939.n0 173.817
R18240 a_8422_1939.n1 a_8422_1939.t1 20.826
R18241 a_8422_1939.n2 a_8422_1939.n1 20.689
R18242 a_13230_n4114.t1 a_13230_n4114.t0 336.812
R18243 RWLB[7].n0 RWLB[7].t0 154.228
R18244 RWLB[7].n14 RWLB[7].t1 149.249
R18245 RWLB[7].n13 RWLB[7].t3 149.249
R18246 RWLB[7].n12 RWLB[7].t14 149.249
R18247 RWLB[7].n11 RWLB[7].t8 149.249
R18248 RWLB[7].n10 RWLB[7].t2 149.249
R18249 RWLB[7].n9 RWLB[7].t5 149.249
R18250 RWLB[7].n8 RWLB[7].t6 149.249
R18251 RWLB[7].n7 RWLB[7].t11 149.249
R18252 RWLB[7].n6 RWLB[7].t4 149.249
R18253 RWLB[7].n5 RWLB[7].t9 149.249
R18254 RWLB[7].n4 RWLB[7].t10 149.249
R18255 RWLB[7].n3 RWLB[7].t15 149.249
R18256 RWLB[7].n2 RWLB[7].t7 149.249
R18257 RWLB[7].n1 RWLB[7].t13 149.249
R18258 RWLB[7].n0 RWLB[7].t12 149.249
R18259 RWLB[7] RWLB[7].n14 47.816
R18260 RWLB[7].n1 RWLB[7].n0 4.979
R18261 RWLB[7].n2 RWLB[7].n1 4.979
R18262 RWLB[7].n3 RWLB[7].n2 4.979
R18263 RWLB[7].n4 RWLB[7].n3 4.979
R18264 RWLB[7].n5 RWLB[7].n4 4.979
R18265 RWLB[7].n6 RWLB[7].n5 4.979
R18266 RWLB[7].n7 RWLB[7].n6 4.979
R18267 RWLB[7].n8 RWLB[7].n7 4.979
R18268 RWLB[7].n9 RWLB[7].n8 4.979
R18269 RWLB[7].n10 RWLB[7].n9 4.979
R18270 RWLB[7].n11 RWLB[7].n10 4.979
R18271 RWLB[7].n12 RWLB[7].n11 4.979
R18272 RWLB[7].n13 RWLB[7].n12 4.979
R18273 RWLB[7].n14 RWLB[7].n13 4.979
R18274 a_8915_n953.t45 a_8915_n953.n46 176.385
R18275 a_8915_n953.n22 a_8915_n953.t7 67.378
R18276 a_8915_n953.n0 a_8915_n953.t4 66.92
R18277 a_8915_n953.n1 a_8915_n953.t11 66.92
R18278 a_8915_n953.n2 a_8915_n953.t16 66.92
R18279 a_8915_n953.n3 a_8915_n953.t8 66.92
R18280 a_8915_n953.n4 a_8915_n953.t0 66.92
R18281 a_8915_n953.n5 a_8915_n953.t21 66.92
R18282 a_8915_n953.n6 a_8915_n953.t48 66.92
R18283 a_8915_n953.n7 a_8915_n953.t31 66.92
R18284 a_8915_n953.n8 a_8915_n953.t23 66.92
R18285 a_8915_n953.n9 a_8915_n953.t37 66.92
R18286 a_8915_n953.n10 a_8915_n953.t35 66.92
R18287 a_8915_n953.n11 a_8915_n953.t19 66.92
R18288 a_8915_n953.n12 a_8915_n953.t32 66.92
R18289 a_8915_n953.n13 a_8915_n953.t36 66.92
R18290 a_8915_n953.n14 a_8915_n953.t34 66.92
R18291 a_8915_n953.n15 a_8915_n953.t25 66.92
R18292 a_8915_n953.n16 a_8915_n953.t17 66.92
R18293 a_8915_n953.n17 a_8915_n953.t28 66.92
R18294 a_8915_n953.n18 a_8915_n953.t26 66.92
R18295 a_8915_n953.n19 a_8915_n953.t29 66.92
R18296 a_8915_n953.n20 a_8915_n953.t2 66.92
R18297 a_8915_n953.n21 a_8915_n953.t14 66.92
R18298 a_8915_n953.n22 a_8915_n953.t5 66.92
R18299 a_8915_n953.n23 a_8915_n953.t15 65.518
R18300 a_8915_n953.n45 a_8915_n953.t1 63.519
R18301 a_8915_n953.n44 a_8915_n953.t9 63.519
R18302 a_8915_n953.n43 a_8915_n953.t3 63.519
R18303 a_8915_n953.n42 a_8915_n953.t13 63.519
R18304 a_8915_n953.n41 a_8915_n953.t43 63.519
R18305 a_8915_n953.n40 a_8915_n953.t40 63.519
R18306 a_8915_n953.n39 a_8915_n953.t24 63.519
R18307 a_8915_n953.n38 a_8915_n953.t42 63.519
R18308 a_8915_n953.n37 a_8915_n953.t20 63.519
R18309 a_8915_n953.n36 a_8915_n953.t27 63.519
R18310 a_8915_n953.n35 a_8915_n953.t39 63.519
R18311 a_8915_n953.n34 a_8915_n953.t46 63.519
R18312 a_8915_n953.n33 a_8915_n953.t38 63.519
R18313 a_8915_n953.n32 a_8915_n953.t22 63.519
R18314 a_8915_n953.n31 a_8915_n953.t18 63.519
R18315 a_8915_n953.n30 a_8915_n953.t47 63.519
R18316 a_8915_n953.n29 a_8915_n953.t44 63.519
R18317 a_8915_n953.n28 a_8915_n953.t41 63.519
R18318 a_8915_n953.n27 a_8915_n953.t33 63.519
R18319 a_8915_n953.n26 a_8915_n953.t30 63.519
R18320 a_8915_n953.n25 a_8915_n953.t10 63.519
R18321 a_8915_n953.n24 a_8915_n953.t6 63.519
R18322 a_8915_n953.n23 a_8915_n953.t12 63.519
R18323 a_8915_n953.n46 a_8915_n953.n45 18.144
R18324 a_8915_n953.n46 a_8915_n953.n0 17.125
R18325 a_8915_n953.n44 a_8915_n953.n43 2.524
R18326 a_8915_n953.n24 a_8915_n953.n23 2.498
R18327 a_8915_n953.n21 a_8915_n953.n22 2.495
R18328 a_8915_n953.n1 a_8915_n953.n2 2.459
R18329 a_8915_n953.n38 a_8915_n953.n37 2.364
R18330 a_8915_n953.n30 a_8915_n953.n29 2.355
R18331 a_8915_n953.n7 a_8915_n953.n8 2.299
R18332 a_8915_n953.n15 a_8915_n953.n16 2.29
R18333 a_8915_n953.n16 a_8915_n953.n17 2.057
R18334 a_8915_n953.n8 a_8915_n953.n9 2.057
R18335 a_8915_n953.n2 a_8915_n953.n3 2.057
R18336 a_8915_n953.n0 a_8915_n953.n1 2.057
R18337 a_8915_n953.n45 a_8915_n953.n44 1.998
R18338 a_8915_n953.n43 a_8915_n953.n42 1.998
R18339 a_8915_n953.n42 a_8915_n953.n41 1.998
R18340 a_8915_n953.n41 a_8915_n953.n40 1.998
R18341 a_8915_n953.n40 a_8915_n953.n39 1.998
R18342 a_8915_n953.n39 a_8915_n953.n38 1.998
R18343 a_8915_n953.n37 a_8915_n953.n36 1.998
R18344 a_8915_n953.n36 a_8915_n953.n35 1.998
R18345 a_8915_n953.n35 a_8915_n953.n34 1.998
R18346 a_8915_n953.n34 a_8915_n953.n33 1.998
R18347 a_8915_n953.n33 a_8915_n953.n32 1.998
R18348 a_8915_n953.n32 a_8915_n953.n31 1.998
R18349 a_8915_n953.n31 a_8915_n953.n30 1.998
R18350 a_8915_n953.n29 a_8915_n953.n28 1.998
R18351 a_8915_n953.n28 a_8915_n953.n27 1.998
R18352 a_8915_n953.n27 a_8915_n953.n26 1.998
R18353 a_8915_n953.n26 a_8915_n953.n25 1.998
R18354 a_8915_n953.n25 a_8915_n953.n24 1.998
R18355 a_8915_n953.n20 a_8915_n953.n21 1.995
R18356 a_8915_n953.n19 a_8915_n953.n20 1.995
R18357 a_8915_n953.n18 a_8915_n953.n19 1.995
R18358 a_8915_n953.n17 a_8915_n953.n18 1.995
R18359 a_8915_n953.n14 a_8915_n953.n15 1.995
R18360 a_8915_n953.n13 a_8915_n953.n14 1.995
R18361 a_8915_n953.n12 a_8915_n953.n13 1.995
R18362 a_8915_n953.n11 a_8915_n953.n12 1.995
R18363 a_8915_n953.n10 a_8915_n953.n11 1.995
R18364 a_8915_n953.n9 a_8915_n953.n10 1.995
R18365 a_8915_n953.n6 a_8915_n953.n7 1.995
R18366 a_8915_n953.n5 a_8915_n953.n6 1.995
R18367 a_8915_n953.n4 a_8915_n953.n5 1.995
R18368 a_8915_n953.n3 a_8915_n953.n4 1.995
R18369 a_9367_1939.t0 a_9367_1939.t1 242.857
R18370 a_4302_437.n0 a_4302_437.t2 362.857
R18371 a_4302_437.t3 a_4302_437.t5 337.399
R18372 a_4302_437.t5 a_4302_437.t4 298.839
R18373 a_4302_437.n0 a_4302_437.t3 280.405
R18374 a_4302_437.n1 a_4302_437.t1 200
R18375 a_4302_437.n1 a_4302_437.n0 172.311
R18376 a_4302_437.n2 a_4302_437.n1 24
R18377 a_4302_437.n1 a_4302_437.t0 21.212
R18378 a_4397_452.n0 a_4397_452.t2 358.166
R18379 a_4397_452.t4 a_4397_452.t3 337.399
R18380 a_4397_452.t3 a_4397_452.t5 285.986
R18381 a_4397_452.n0 a_4397_452.t4 282.573
R18382 a_4397_452.n1 a_4397_452.t0 202.857
R18383 a_4397_452.n1 a_4397_452.n0 173.817
R18384 a_4397_452.n1 a_4397_452.t1 20.826
R18385 a_4397_452.n2 a_4397_452.n1 20.689
R18386 a_7190_n812.t0 a_7190_n812.t1 242.857
R18387 a_2097_3666.n0 a_2097_3666.t1 358.166
R18388 a_2097_3666.t4 a_2097_3666.t5 337.399
R18389 a_2097_3666.t5 a_2097_3666.t3 285.986
R18390 a_2097_3666.n0 a_2097_3666.t4 282.573
R18391 a_2097_3666.n1 a_2097_3666.t2 202.857
R18392 a_2097_3666.n1 a_2097_3666.n0 173.817
R18393 a_2097_3666.n1 a_2097_3666.t0 20.826
R18394 a_2097_3666.n2 a_2097_3666.n1 20.689
R18395 a_2467_3666.t0 a_2467_3666.t1 242.857
R18396 RWLB[15].n0 RWLB[15].t14 154.228
R18397 RWLB[15].n14 RWLB[15].t3 149.249
R18398 RWLB[15].n13 RWLB[15].t2 149.249
R18399 RWLB[15].n12 RWLB[15].t10 149.249
R18400 RWLB[15].n11 RWLB[15].t6 149.249
R18401 RWLB[15].n10 RWLB[15].t13 149.249
R18402 RWLB[15].n9 RWLB[15].t12 149.249
R18403 RWLB[15].n8 RWLB[15].t0 149.249
R18404 RWLB[15].n7 RWLB[15].t15 149.249
R18405 RWLB[15].n6 RWLB[15].t8 149.249
R18406 RWLB[15].n5 RWLB[15].t7 149.249
R18407 RWLB[15].n4 RWLB[15].t9 149.249
R18408 RWLB[15].n3 RWLB[15].t4 149.249
R18409 RWLB[15].n2 RWLB[15].t1 149.249
R18410 RWLB[15].n1 RWLB[15].t11 149.249
R18411 RWLB[15].n0 RWLB[15].t5 149.249
R18412 RWLB[15] RWLB[15].n14 47.816
R18413 RWLB[15].n1 RWLB[15].n0 4.979
R18414 RWLB[15].n2 RWLB[15].n1 4.979
R18415 RWLB[15].n3 RWLB[15].n2 4.979
R18416 RWLB[15].n4 RWLB[15].n3 4.979
R18417 RWLB[15].n5 RWLB[15].n4 4.979
R18418 RWLB[15].n6 RWLB[15].n5 4.979
R18419 RWLB[15].n7 RWLB[15].n6 4.979
R18420 RWLB[15].n8 RWLB[15].n7 4.979
R18421 RWLB[15].n9 RWLB[15].n8 4.979
R18422 RWLB[15].n10 RWLB[15].n9 4.979
R18423 RWLB[15].n11 RWLB[15].n10 4.979
R18424 RWLB[15].n12 RWLB[15].n11 4.979
R18425 RWLB[15].n13 RWLB[15].n12 4.979
R18426 RWLB[15].n14 RWLB[15].n13 4.979
R18427 a_4192_n30.t0 a_4192_n30.t1 242.857
R18428 a_4877_3169.n0 a_4877_3169.t2 362.857
R18429 a_4877_3169.t5 a_4877_3169.t4 337.399
R18430 a_4877_3169.t4 a_4877_3169.t3 298.839
R18431 a_4877_3169.n0 a_4877_3169.t5 280.405
R18432 a_4877_3169.n1 a_4877_3169.t0 200
R18433 a_4877_3169.n1 a_4877_3169.n0 172.311
R18434 a_4877_3169.n2 a_4877_3169.n1 24
R18435 a_4877_3169.n1 a_4877_3169.t1 21.212
R18436 a_4890_3184.t0 a_4890_3184.t1 242.857
R18437 a_3420_4887.n25 a_3420_4887.t27 561.971
R18438 a_3420_4887.n0 a_3420_4887.t5 449.944
R18439 a_3420_4887.t14 a_3420_4887.n25 108.636
R18440 a_3420_4887.n0 a_3420_4887.t6 74.821
R18441 a_3420_4887.n24 a_3420_4887.t20 63.519
R18442 a_3420_4887.n23 a_3420_4887.t1 63.519
R18443 a_3420_4887.n22 a_3420_4887.t13 63.519
R18444 a_3420_4887.n21 a_3420_4887.t15 63.519
R18445 a_3420_4887.n20 a_3420_4887.t22 63.519
R18446 a_3420_4887.n19 a_3420_4887.t18 63.519
R18447 a_3420_4887.n18 a_3420_4887.t19 63.519
R18448 a_3420_4887.n17 a_3420_4887.t10 63.519
R18449 a_3420_4887.n16 a_3420_4887.t4 63.519
R18450 a_3420_4887.n15 a_3420_4887.t8 63.519
R18451 a_3420_4887.n14 a_3420_4887.t21 63.519
R18452 a_3420_4887.n13 a_3420_4887.t23 63.519
R18453 a_3420_4887.n12 a_3420_4887.t17 63.519
R18454 a_3420_4887.n11 a_3420_4887.t11 63.519
R18455 a_3420_4887.n10 a_3420_4887.t12 63.519
R18456 a_3420_4887.n9 a_3420_4887.t24 63.519
R18457 a_3420_4887.n8 a_3420_4887.t0 63.519
R18458 a_3420_4887.n7 a_3420_4887.t3 63.519
R18459 a_3420_4887.n6 a_3420_4887.t2 63.519
R18460 a_3420_4887.n5 a_3420_4887.t26 63.519
R18461 a_3420_4887.n4 a_3420_4887.t9 63.519
R18462 a_3420_4887.n3 a_3420_4887.t16 63.519
R18463 a_3420_4887.n2 a_3420_4887.t25 63.519
R18464 a_3420_4887.n1 a_3420_4887.t7 63.519
R18465 a_3420_4887.n1 a_3420_4887.n0 8.619
R18466 a_3420_4887.n25 a_3420_4887.n24 2.946
R18467 a_3420_4887.n23 a_3420_4887.n22 2.524
R18468 a_3420_4887.n3 a_3420_4887.n2 2.498
R18469 a_3420_4887.n17 a_3420_4887.n16 2.364
R18470 a_3420_4887.n9 a_3420_4887.n8 2.355
R18471 a_3420_4887.n24 a_3420_4887.n23 1.998
R18472 a_3420_4887.n22 a_3420_4887.n21 1.998
R18473 a_3420_4887.n21 a_3420_4887.n20 1.998
R18474 a_3420_4887.n20 a_3420_4887.n19 1.998
R18475 a_3420_4887.n19 a_3420_4887.n18 1.998
R18476 a_3420_4887.n18 a_3420_4887.n17 1.998
R18477 a_3420_4887.n16 a_3420_4887.n15 1.998
R18478 a_3420_4887.n15 a_3420_4887.n14 1.998
R18479 a_3420_4887.n14 a_3420_4887.n13 1.998
R18480 a_3420_4887.n13 a_3420_4887.n12 1.998
R18481 a_3420_4887.n12 a_3420_4887.n11 1.998
R18482 a_3420_4887.n11 a_3420_4887.n10 1.998
R18483 a_3420_4887.n10 a_3420_4887.n9 1.998
R18484 a_3420_4887.n8 a_3420_4887.n7 1.998
R18485 a_3420_4887.n7 a_3420_4887.n6 1.998
R18486 a_3420_4887.n6 a_3420_4887.n5 1.998
R18487 a_3420_4887.n5 a_3420_4887.n4 1.998
R18488 a_3420_4887.n4 a_3420_4887.n3 1.998
R18489 a_3420_4887.n2 a_3420_4887.n1 1.998
R18490 a_3152_1924.n0 a_3152_1924.t0 362.857
R18491 a_3152_1924.t3 a_3152_1924.t4 337.399
R18492 a_3152_1924.t4 a_3152_1924.t5 298.839
R18493 a_3152_1924.n0 a_3152_1924.t3 280.405
R18494 a_3152_1924.n1 a_3152_1924.t2 200
R18495 a_3152_1924.n1 a_3152_1924.n0 172.311
R18496 a_3152_1924.n2 a_3152_1924.n1 24
R18497 a_3152_1924.n1 a_3152_1924.t1 21.212
R18498 WWL[15].n0 WWL[15].t2 262.032
R18499 WWL[15].n29 WWL[15].t14 260.715
R18500 WWL[15].n27 WWL[15].t12 260.715
R18501 WWL[15].n25 WWL[15].t5 260.715
R18502 WWL[15].n23 WWL[15].t18 260.715
R18503 WWL[15].n21 WWL[15].t13 260.715
R18504 WWL[15].n19 WWL[15].t31 260.715
R18505 WWL[15].n17 WWL[15].t19 260.715
R18506 WWL[15].n15 WWL[15].t3 260.715
R18507 WWL[15].n13 WWL[15].t23 260.715
R18508 WWL[15].n11 WWL[15].t21 260.715
R18509 WWL[15].n9 WWL[15].t4 260.715
R18510 WWL[15].n7 WWL[15].t24 260.715
R18511 WWL[15].n5 WWL[15].t11 260.715
R18512 WWL[15].n3 WWL[15].t30 260.715
R18513 WWL[15].n1 WWL[15].t26 260.715
R18514 WWL[15].n30 WWL[15].t10 259.254
R18515 WWL[15].n28 WWL[15].t0 259.254
R18516 WWL[15].n26 WWL[15].t8 259.254
R18517 WWL[15].n24 WWL[15].t9 259.254
R18518 WWL[15].n22 WWL[15].t20 259.254
R18519 WWL[15].n20 WWL[15].t22 259.254
R18520 WWL[15].n18 WWL[15].t28 259.254
R18521 WWL[15].n16 WWL[15].t29 259.254
R18522 WWL[15].n14 WWL[15].t6 259.254
R18523 WWL[15].n12 WWL[15].t7 259.254
R18524 WWL[15].n10 WWL[15].t25 259.254
R18525 WWL[15].n8 WWL[15].t17 259.254
R18526 WWL[15].n6 WWL[15].t1 259.254
R18527 WWL[15].n4 WWL[15].t27 259.254
R18528 WWL[15].n2 WWL[15].t15 259.254
R18529 WWL[15].n0 WWL[15].t16 259.254
R18530 WWL[15] WWL[15].n30 44.647
R18531 WWL[15].n1 WWL[15].n0 3.576
R18532 WWL[15].n3 WWL[15].n2 3.576
R18533 WWL[15].n5 WWL[15].n4 3.576
R18534 WWL[15].n7 WWL[15].n6 3.576
R18535 WWL[15].n9 WWL[15].n8 3.576
R18536 WWL[15].n11 WWL[15].n10 3.576
R18537 WWL[15].n13 WWL[15].n12 3.576
R18538 WWL[15].n15 WWL[15].n14 3.576
R18539 WWL[15].n17 WWL[15].n16 3.576
R18540 WWL[15].n19 WWL[15].n18 3.576
R18541 WWL[15].n21 WWL[15].n20 3.576
R18542 WWL[15].n23 WWL[15].n22 3.576
R18543 WWL[15].n25 WWL[15].n24 3.576
R18544 WWL[15].n27 WWL[15].n26 3.576
R18545 WWL[15].n29 WWL[15].n28 3.576
R18546 WWL[15].n2 WWL[15].n1 1.317
R18547 WWL[15].n4 WWL[15].n3 1.317
R18548 WWL[15].n6 WWL[15].n5 1.317
R18549 WWL[15].n8 WWL[15].n7 1.317
R18550 WWL[15].n10 WWL[15].n9 1.317
R18551 WWL[15].n12 WWL[15].n11 1.317
R18552 WWL[15].n14 WWL[15].n13 1.317
R18553 WWL[15].n16 WWL[15].n15 1.317
R18554 WWL[15].n18 WWL[15].n17 1.317
R18555 WWL[15].n20 WWL[15].n19 1.317
R18556 WWL[15].n22 WWL[15].n21 1.317
R18557 WWL[15].n24 WWL[15].n23 1.317
R18558 WWL[15].n26 WWL[15].n25 1.317
R18559 WWL[15].n28 WWL[15].n27 1.317
R18560 WWL[15].n30 WWL[15].n29 1.317
R18561 a_947_n30.n0 a_947_n30.t2 358.166
R18562 a_947_n30.t5 a_947_n30.t4 337.399
R18563 a_947_n30.t4 a_947_n30.t3 285.986
R18564 a_947_n30.n0 a_947_n30.t5 282.573
R18565 a_947_n30.n1 a_947_n30.t0 202.857
R18566 a_947_n30.n1 a_947_n30.n0 173.817
R18567 a_947_n30.n1 a_947_n30.t1 20.826
R18568 a_947_n30.n2 a_947_n30.n1 20.689
R18569 a_2097_n512.n0 a_2097_n512.t1 358.166
R18570 a_2097_n512.t5 a_2097_n512.t3 337.399
R18571 a_2097_n512.t3 a_2097_n512.t4 285.986
R18572 a_2097_n512.n0 a_2097_n512.t5 282.573
R18573 a_2097_n512.n1 a_2097_n512.t0 202.857
R18574 a_2097_n512.n1 a_2097_n512.n0 173.817
R18575 a_2097_n512.n1 a_2097_n512.t2 20.826
R18576 a_2097_n512.n2 a_2097_n512.n1 20.689
R18577 a_2002_n527.n0 a_2002_n527.t1 362.857
R18578 a_2002_n527.t3 a_2002_n527.t5 337.399
R18579 a_2002_n527.t5 a_2002_n527.t4 298.839
R18580 a_2002_n527.n0 a_2002_n527.t3 280.405
R18581 a_2002_n527.n1 a_2002_n527.t2 200
R18582 a_2002_n527.n1 a_2002_n527.n0 172.311
R18583 a_2002_n527.n2 a_2002_n527.n1 24
R18584 a_2002_n527.n1 a_2002_n527.t0 21.212
R18585 a_2590_4686.t0 a_2590_4686.t1 242.857
R18586 a_852_4133.n0 a_852_4133.t1 362.857
R18587 a_852_4133.t3 a_852_4133.t4 337.399
R18588 a_852_4133.t4 a_852_4133.t5 298.839
R18589 a_852_4133.n0 a_852_4133.t3 280.405
R18590 a_852_4133.n1 a_852_4133.t0 200
R18591 a_852_4133.n1 a_852_4133.n0 172.311
R18592 a_852_4133.n2 a_852_4133.n1 24
R18593 a_852_4133.n1 a_852_4133.t2 21.212
R18594 a_947_4148.n0 a_947_4148.t1 358.166
R18595 a_947_4148.t4 a_947_4148.t5 337.399
R18596 a_947_4148.t5 a_947_4148.t3 285.986
R18597 a_947_4148.n0 a_947_4148.t4 282.573
R18598 a_947_4148.n1 a_947_4148.t2 202.857
R18599 a_947_4148.n1 a_947_4148.n0 173.817
R18600 a_947_4148.n1 a_947_4148.t0 20.826
R18601 a_947_4148.n2 a_947_4148.n1 20.689
R18602 a_7177_3169.n0 a_7177_3169.t1 362.857
R18603 a_7177_3169.t3 a_7177_3169.t4 337.399
R18604 a_7177_3169.t4 a_7177_3169.t5 298.839
R18605 a_7177_3169.n0 a_7177_3169.t3 280.405
R18606 a_7177_3169.n1 a_7177_3169.t0 200
R18607 a_7177_3169.n1 a_7177_3169.n0 172.311
R18608 a_7177_3169.n2 a_7177_3169.n1 24
R18609 a_7177_3169.n1 a_7177_3169.t2 21.212
R18610 a_7272_3184.n0 a_7272_3184.t2 358.166
R18611 a_7272_3184.t4 a_7272_3184.t3 337.399
R18612 a_7272_3184.t3 a_7272_3184.t5 285.986
R18613 a_7272_3184.n0 a_7272_3184.t4 282.573
R18614 a_7272_3184.n1 a_7272_3184.t0 202.857
R18615 a_7272_3184.n1 a_7272_3184.n0 173.817
R18616 a_7272_3184.n1 a_7272_3184.t1 20.826
R18617 a_7272_3184.n2 a_7272_3184.n1 20.689
R18618 a_310_n1371.n1 a_310_n1371.t3 550.94
R18619 a_310_n1371.n1 a_310_n1371.t4 500.621
R18620 a_310_n1371.t1 a_310_n1371.n2 192.787
R18621 a_310_n1371.n0 a_310_n1371.t0 163.997
R18622 a_310_n1371.n2 a_310_n1371.n1 149.035
R18623 a_310_n1371.n0 a_310_n1371.t2 54.068
R18624 a_310_n1371.n2 a_310_n1371.n0 17.317
R18625 a_3822_1698.n0 a_3822_1698.t1 358.166
R18626 a_3822_1698.t4 a_3822_1698.t3 337.399
R18627 a_3822_1698.t3 a_3822_1698.t5 285.986
R18628 a_3822_1698.n0 a_3822_1698.t4 282.573
R18629 a_3822_1698.n1 a_3822_1698.t0 202.857
R18630 a_3822_1698.n1 a_3822_1698.n0 173.817
R18631 a_3822_1698.n1 a_3822_1698.t2 20.826
R18632 a_3822_1698.n2 a_3822_1698.n1 20.689
R18633 a_3727_1683.n0 a_3727_1683.t2 362.857
R18634 a_3727_1683.t3 a_3727_1683.t4 337.399
R18635 a_3727_1683.t4 a_3727_1683.t5 298.839
R18636 a_3727_1683.n0 a_3727_1683.t3 280.405
R18637 a_3727_1683.n1 a_3727_1683.t0 200
R18638 a_3727_1683.n1 a_3727_1683.n0 172.311
R18639 a_3727_1683.n2 a_3727_1683.n1 24
R18640 a_3727_1683.n1 a_3727_1683.t1 21.212
R18641 a_3247_1216.n0 a_3247_1216.t2 358.166
R18642 a_3247_1216.t5 a_3247_1216.t3 337.399
R18643 a_3247_1216.t3 a_3247_1216.t4 285.986
R18644 a_3247_1216.n0 a_3247_1216.t5 282.573
R18645 a_3247_1216.n1 a_3247_1216.t1 202.857
R18646 a_3247_1216.n1 a_3247_1216.n0 173.817
R18647 a_3247_1216.n1 a_3247_1216.t0 20.826
R18648 a_3247_1216.n2 a_3247_1216.n1 20.689
R18649 a_3152_1201.n0 a_3152_1201.t2 362.857
R18650 a_3152_1201.t3 a_3152_1201.t4 337.399
R18651 a_3152_1201.t4 a_3152_1201.t5 298.839
R18652 a_3152_1201.n0 a_3152_1201.t3 280.405
R18653 a_3152_1201.n1 a_3152_1201.t0 200
R18654 a_3152_1201.n1 a_3152_1201.n0 172.311
R18655 a_3152_1201.n2 a_3152_1201.n1 24
R18656 a_3152_1201.n1 a_3152_1201.t1 21.212
R18657 ADC6_OUT[3].n0 ADC6_OUT[3].t3 1355.37
R18658 ADC6_OUT[3].n0 ADC6_OUT[3].t4 820.859
R18659 ADC6_OUT[3].n3 ADC6_OUT[3].t0 336.667
R18660 ADC6_OUT[3].n2 ADC6_OUT[3].t2 266.644
R18661 ADC6_OUT[3].n1 ADC6_OUT[3].n0 149.035
R18662 ADC6_OUT[3].n3 ADC6_OUT[3].n2 47.435
R18663 ADC6_OUT[3].n1 ADC6_OUT[3].t1 45.968
R18664 ADC6_OUT[3] ADC6_OUT[3].n3 22.213
R18665 ADC6_OUT[3].n2 ADC6_OUT[3].n1 17.317
R18666 a_4952_n2234.n2 a_4952_n2234.t1 282.97
R18667 a_4952_n2234.n1 a_4952_n2234.t3 240.683
R18668 a_4952_n2234.n0 a_4952_n2234.t4 209.208
R18669 a_4952_n2234.n0 a_4952_n2234.t2 194.167
R18670 a_4952_n2234.t0 a_4952_n2234.n2 183.404
R18671 a_4952_n2234.n1 a_4952_n2234.n0 14.805
R18672 a_4952_n2234.n2 a_4952_n2234.n1 6.415
R18673 a_5075_n2132.n0 a_5075_n2132.t2 489.336
R18674 a_5075_n2132.n0 a_5075_n2132.t1 243.258
R18675 a_5075_n2132.t0 a_5075_n2132.n0 214.415
R18676 a_2002_960.n0 a_2002_960.t2 362.857
R18677 a_2002_960.t4 a_2002_960.t3 337.399
R18678 a_2002_960.t3 a_2002_960.t5 298.839
R18679 a_2002_960.n0 a_2002_960.t4 280.405
R18680 a_2002_960.n1 a_2002_960.t0 200
R18681 a_2002_960.n1 a_2002_960.n0 172.311
R18682 a_2002_960.n2 a_2002_960.n1 24
R18683 a_2002_960.n1 a_2002_960.t1 21.212
R18684 a_2097_975.n0 a_2097_975.t1 358.166
R18685 a_2097_975.t4 a_2097_975.t5 337.399
R18686 a_2097_975.t5 a_2097_975.t3 285.986
R18687 a_2097_975.n0 a_2097_975.t4 282.573
R18688 a_2097_975.n1 a_2097_975.t2 202.857
R18689 a_2097_975.n1 a_2097_975.n0 173.817
R18690 a_2097_975.n1 a_2097_975.t0 20.826
R18691 a_2097_975.n2 a_2097_975.n1 20.689
R18692 a_1522_n271.n0 a_1522_n271.t1 358.166
R18693 a_1522_n271.t5 a_1522_n271.t4 337.399
R18694 a_1522_n271.t4 a_1522_n271.t3 285.986
R18695 a_1522_n271.n0 a_1522_n271.t5 282.573
R18696 a_1522_n271.n1 a_1522_n271.t0 202.857
R18697 a_1522_n271.n1 a_1522_n271.n0 173.817
R18698 a_1522_n271.n1 a_1522_n271.t2 20.826
R18699 a_1522_n271.n2 a_1522_n271.n1 20.689
R18700 a_1892_n271.t0 a_1892_n271.t1 242.857
R18701 a_1427_n827.n0 a_1427_n827.t1 362.857
R18702 a_1427_n827.t4 a_1427_n827.t5 337.399
R18703 a_1427_n827.t5 a_1427_n827.t3 298.839
R18704 a_1427_n827.n0 a_1427_n827.t4 280.405
R18705 a_1427_n827.n1 a_1427_n827.t0 200
R18706 a_1427_n827.n1 a_1427_n827.n0 172.311
R18707 a_1427_n827.n2 a_1427_n827.n1 24
R18708 a_1427_n827.n1 a_1427_n827.t2 21.212
R18709 a_1440_n812.t0 a_1440_n812.t1 242.857
R18710 a_2002_2406.n0 a_2002_2406.t1 362.857
R18711 a_2002_2406.t3 a_2002_2406.t5 337.399
R18712 a_2002_2406.t5 a_2002_2406.t4 298.839
R18713 a_2002_2406.n0 a_2002_2406.t3 280.405
R18714 a_2002_2406.n1 a_2002_2406.t0 200
R18715 a_2002_2406.n1 a_2002_2406.n0 172.311
R18716 a_2002_2406.n2 a_2002_2406.n1 24
R18717 a_2002_2406.n1 a_2002_2406.t2 21.212
R18718 a_2097_2421.n0 a_2097_2421.t1 358.166
R18719 a_2097_2421.t5 a_2097_2421.t3 337.399
R18720 a_2097_2421.t3 a_2097_2421.t4 285.986
R18721 a_2097_2421.n0 a_2097_2421.t5 282.573
R18722 a_2097_2421.n1 a_2097_2421.t2 202.857
R18723 a_2097_2421.n1 a_2097_2421.n0 173.817
R18724 a_2097_2421.n1 a_2097_2421.t0 20.826
R18725 a_2097_2421.n2 a_2097_2421.n1 20.689
R18726 WWL[8].n0 WWL[8].t14 262.032
R18727 WWL[8].n29 WWL[8].t17 260.715
R18728 WWL[8].n27 WWL[8].t20 260.715
R18729 WWL[8].n25 WWL[8].t2 260.715
R18730 WWL[8].n23 WWL[8].t28 260.715
R18731 WWL[8].n21 WWL[8].t8 260.715
R18732 WWL[8].n19 WWL[8].t25 260.715
R18733 WWL[8].n17 WWL[8].t16 260.715
R18734 WWL[8].n15 WWL[8].t31 260.715
R18735 WWL[8].n13 WWL[8].t21 260.715
R18736 WWL[8].n11 WWL[8].t29 260.715
R18737 WWL[8].n9 WWL[8].t18 260.715
R18738 WWL[8].n7 WWL[8].t0 260.715
R18739 WWL[8].n5 WWL[8].t26 260.715
R18740 WWL[8].n3 WWL[8].t9 260.715
R18741 WWL[8].n1 WWL[8].t22 260.715
R18742 WWL[8].n30 WWL[8].t1 259.254
R18743 WWL[8].n28 WWL[8].t7 259.254
R18744 WWL[8].n26 WWL[8].t19 259.254
R18745 WWL[8].n24 WWL[8].t3 259.254
R18746 WWL[8].n22 WWL[8].t27 259.254
R18747 WWL[8].n20 WWL[8].t10 259.254
R18748 WWL[8].n18 WWL[8].t23 259.254
R18749 WWL[8].n16 WWL[8].t5 259.254
R18750 WWL[8].n14 WWL[8].t30 259.254
R18751 WWL[8].n12 WWL[8].t13 259.254
R18752 WWL[8].n10 WWL[8].t4 259.254
R18753 WWL[8].n8 WWL[8].t11 259.254
R18754 WWL[8].n6 WWL[8].t12 259.254
R18755 WWL[8].n4 WWL[8].t15 259.254
R18756 WWL[8].n2 WWL[8].t6 259.254
R18757 WWL[8].n0 WWL[8].t24 259.254
R18758 WWL[8] WWL[8].n30 44.647
R18759 WWL[8].n1 WWL[8].n0 3.576
R18760 WWL[8].n3 WWL[8].n2 3.576
R18761 WWL[8].n5 WWL[8].n4 3.576
R18762 WWL[8].n7 WWL[8].n6 3.576
R18763 WWL[8].n9 WWL[8].n8 3.576
R18764 WWL[8].n11 WWL[8].n10 3.576
R18765 WWL[8].n13 WWL[8].n12 3.576
R18766 WWL[8].n15 WWL[8].n14 3.576
R18767 WWL[8].n17 WWL[8].n16 3.576
R18768 WWL[8].n19 WWL[8].n18 3.576
R18769 WWL[8].n21 WWL[8].n20 3.576
R18770 WWL[8].n23 WWL[8].n22 3.576
R18771 WWL[8].n25 WWL[8].n24 3.576
R18772 WWL[8].n27 WWL[8].n26 3.576
R18773 WWL[8].n29 WWL[8].n28 3.576
R18774 WWL[8].n2 WWL[8].n1 1.317
R18775 WWL[8].n4 WWL[8].n3 1.317
R18776 WWL[8].n6 WWL[8].n5 1.317
R18777 WWL[8].n8 WWL[8].n7 1.317
R18778 WWL[8].n10 WWL[8].n9 1.317
R18779 WWL[8].n12 WWL[8].n11 1.317
R18780 WWL[8].n14 WWL[8].n13 1.317
R18781 WWL[8].n16 WWL[8].n15 1.317
R18782 WWL[8].n18 WWL[8].n17 1.317
R18783 WWL[8].n20 WWL[8].n19 1.317
R18784 WWL[8].n22 WWL[8].n21 1.317
R18785 WWL[8].n24 WWL[8].n23 1.317
R18786 WWL[8].n26 WWL[8].n25 1.317
R18787 WWL[8].n28 WWL[8].n27 1.317
R18788 WWL[8].n30 WWL[8].n29 1.317
R18789 a_6602_1683.n0 a_6602_1683.t0 362.857
R18790 a_6602_1683.t3 a_6602_1683.t5 337.399
R18791 a_6602_1683.t5 a_6602_1683.t4 298.839
R18792 a_6602_1683.n0 a_6602_1683.t3 280.405
R18793 a_6602_1683.n1 a_6602_1683.t2 200
R18794 a_6602_1683.n1 a_6602_1683.n0 172.311
R18795 a_6602_1683.n2 a_6602_1683.n1 24
R18796 a_6602_1683.n1 a_6602_1683.t1 21.212
R18797 RWL[15].n0 RWL[15].t9 154.243
R18798 RWL[15].n14 RWL[15].t14 149.249
R18799 RWL[15].n13 RWL[15].t7 149.249
R18800 RWL[15].n12 RWL[15].t12 149.249
R18801 RWL[15].n11 RWL[15].t13 149.249
R18802 RWL[15].n10 RWL[15].t1 149.249
R18803 RWL[15].n9 RWL[15].t2 149.249
R18804 RWL[15].n8 RWL[15].t5 149.249
R18805 RWL[15].n7 RWL[15].t6 149.249
R18806 RWL[15].n6 RWL[15].t10 149.249
R18807 RWL[15].n5 RWL[15].t11 149.249
R18808 RWL[15].n4 RWL[15].t3 149.249
R18809 RWL[15].n3 RWL[15].t0 149.249
R18810 RWL[15].n2 RWL[15].t8 149.249
R18811 RWL[15].n1 RWL[15].t4 149.249
R18812 RWL[15].n0 RWL[15].t15 149.249
R18813 RWL[15] RWL[15].n14 42.872
R18814 RWL[15].n1 RWL[15].n0 4.994
R18815 RWL[15].n2 RWL[15].n1 4.994
R18816 RWL[15].n3 RWL[15].n2 4.994
R18817 RWL[15].n4 RWL[15].n3 4.994
R18818 RWL[15].n5 RWL[15].n4 4.994
R18819 RWL[15].n6 RWL[15].n5 4.994
R18820 RWL[15].n7 RWL[15].n6 4.994
R18821 RWL[15].n8 RWL[15].n7 4.994
R18822 RWL[15].n9 RWL[15].n8 4.994
R18823 RWL[15].n10 RWL[15].n9 4.994
R18824 RWL[15].n11 RWL[15].n10 4.994
R18825 RWL[15].n12 RWL[15].n11 4.994
R18826 RWL[15].n13 RWL[15].n12 4.994
R18827 RWL[15].n14 RWL[15].n13 4.994
R18828 a_6615_n30.t0 a_6615_n30.t1 242.857
R18829 a_8915_n512.t0 a_8915_n512.t1 242.857
R18830 a_5452_3651.n0 a_5452_3651.t0 362.857
R18831 a_5452_3651.t3 a_5452_3651.t4 337.399
R18832 a_5452_3651.t4 a_5452_3651.t5 298.839
R18833 a_5452_3651.n0 a_5452_3651.t3 280.405
R18834 a_5452_3651.n1 a_5452_3651.t2 200
R18835 a_5452_3651.n1 a_5452_3651.n0 172.311
R18836 a_5452_3651.n2 a_5452_3651.n1 24
R18837 a_5452_3651.n1 a_5452_3651.t1 21.212
R18838 a_2178_n2086.t0 a_2178_n2086.t1 34.8
R18839 a_3165_4445.t0 a_3165_4445.t1 242.857
R18840 a_6027_4430.n0 a_6027_4430.t1 362.857
R18841 a_6027_4430.t5 a_6027_4430.t3 337.399
R18842 a_6027_4430.t3 a_6027_4430.t4 298.839
R18843 a_6027_4430.n0 a_6027_4430.t5 280.405
R18844 a_6027_4430.n1 a_6027_4430.t2 200
R18845 a_6027_4430.n1 a_6027_4430.n0 172.311
R18846 a_6027_4430.n2 a_6027_4430.n1 24
R18847 a_6027_4430.n1 a_6027_4430.t0 21.212
R18848 a_6122_4445.n0 a_6122_4445.t1 358.166
R18849 a_6122_4445.t4 a_6122_4445.t3 337.399
R18850 a_6122_4445.t3 a_6122_4445.t5 285.986
R18851 a_6122_4445.n0 a_6122_4445.t4 282.573
R18852 a_6122_4445.n1 a_6122_4445.t2 202.857
R18853 a_6122_4445.n1 a_6122_4445.n0 173.817
R18854 a_6122_4445.n1 a_6122_4445.t0 20.826
R18855 a_6122_4445.n2 a_6122_4445.n1 20.689
R18856 RWLB[0].n0 RWLB[0].t15 154.228
R18857 RWLB[0].n14 RWLB[0].t0 149.249
R18858 RWLB[0].n13 RWLB[0].t2 149.249
R18859 RWLB[0].n12 RWLB[0].t13 149.249
R18860 RWLB[0].n11 RWLB[0].t7 149.249
R18861 RWLB[0].n10 RWLB[0].t1 149.249
R18862 RWLB[0].n9 RWLB[0].t4 149.249
R18863 RWLB[0].n8 RWLB[0].t5 149.249
R18864 RWLB[0].n7 RWLB[0].t10 149.249
R18865 RWLB[0].n6 RWLB[0].t3 149.249
R18866 RWLB[0].n5 RWLB[0].t8 149.249
R18867 RWLB[0].n4 RWLB[0].t9 149.249
R18868 RWLB[0].n3 RWLB[0].t14 149.249
R18869 RWLB[0].n2 RWLB[0].t6 149.249
R18870 RWLB[0].n1 RWLB[0].t12 149.249
R18871 RWLB[0].n0 RWLB[0].t11 149.249
R18872 RWLB[0] RWLB[0].n14 47.816
R18873 RWLB[0].n1 RWLB[0].n0 4.979
R18874 RWLB[0].n2 RWLB[0].n1 4.979
R18875 RWLB[0].n3 RWLB[0].n2 4.979
R18876 RWLB[0].n4 RWLB[0].n3 4.979
R18877 RWLB[0].n5 RWLB[0].n4 4.979
R18878 RWLB[0].n6 RWLB[0].n5 4.979
R18879 RWLB[0].n7 RWLB[0].n6 4.979
R18880 RWLB[0].n8 RWLB[0].n7 4.979
R18881 RWLB[0].n9 RWLB[0].n8 4.979
R18882 RWLB[0].n10 RWLB[0].n9 4.979
R18883 RWLB[0].n11 RWLB[0].n10 4.979
R18884 RWLB[0].n12 RWLB[0].n11 4.979
R18885 RWLB[0].n13 RWLB[0].n12 4.979
R18886 RWLB[0].n14 RWLB[0].n13 4.979
R18887 a_742_3666.t0 a_742_3666.t1 242.857
R18888 a_2002_n286.n0 a_2002_n286.t1 362.857
R18889 a_2002_n286.t3 a_2002_n286.t5 337.399
R18890 a_2002_n286.t5 a_2002_n286.t4 298.839
R18891 a_2002_n286.n0 a_2002_n286.t3 280.405
R18892 a_2002_n286.n1 a_2002_n286.t0 200
R18893 a_2002_n286.n1 a_2002_n286.n0 172.311
R18894 a_2002_n286.n2 a_2002_n286.n1 24
R18895 a_2002_n286.n1 a_2002_n286.t2 21.212
R18896 a_2097_n271.n0 a_2097_n271.t1 358.166
R18897 a_2097_n271.t4 a_2097_n271.t5 337.399
R18898 a_2097_n271.t5 a_2097_n271.t3 285.986
R18899 a_2097_n271.n0 a_2097_n271.t4 282.573
R18900 a_2097_n271.n1 a_2097_n271.t2 202.857
R18901 a_2097_n271.n1 a_2097_n271.n0 173.817
R18902 a_2097_n271.n1 a_2097_n271.t0 20.826
R18903 a_2097_n271.n2 a_2097_n271.n1 20.689
R18904 a_n52_n5850.n0 a_n52_n5850.t4 1465.51
R18905 a_n52_n5850.n0 a_n52_n5850.t3 712.44
R18906 a_n52_n5850.n1 a_n52_n5850.t0 375.067
R18907 a_n52_n5850.n1 a_n52_n5850.t1 272.668
R18908 a_n52_n5850.n2 a_n52_n5850.n0 143.764
R18909 a_n52_n5850.t2 a_n52_n5850.n2 78.193
R18910 a_n52_n5850.n2 a_n52_n5850.n1 4.517
R18911 a_277_n1068.n0 a_277_n1068.t1 362.857
R18912 a_277_n1068.t3 a_277_n1068.t4 337.399
R18913 a_277_n1068.t4 a_277_n1068.t5 298.839
R18914 a_277_n1068.n0 a_277_n1068.t3 280.405
R18915 a_277_n1068.n1 a_277_n1068.t2 200
R18916 a_277_n1068.n1 a_277_n1068.n0 172.311
R18917 a_277_n1068.n2 a_277_n1068.n1 24
R18918 a_277_n1068.n1 a_277_n1068.t0 21.212
R18919 a_372_n1053.n0 a_372_n1053.t1 358.166
R18920 a_372_n1053.t5 a_372_n1053.t4 337.399
R18921 a_372_n1053.t4 a_372_n1053.t3 285.986
R18922 a_372_n1053.n0 a_372_n1053.t5 282.573
R18923 a_372_n1053.n1 a_372_n1053.t2 202.857
R18924 a_372_n1053.n1 a_372_n1053.n0 173.817
R18925 a_372_n1053.n1 a_372_n1053.t0 20.826
R18926 a_372_n1053.n2 a_372_n1053.n1 20.689
R18927 a_1522_3425.n0 a_1522_3425.t2 358.166
R18928 a_1522_3425.t5 a_1522_3425.t4 337.399
R18929 a_1522_3425.t4 a_1522_3425.t3 285.986
R18930 a_1522_3425.n0 a_1522_3425.t5 282.573
R18931 a_1522_3425.n1 a_1522_3425.t0 202.857
R18932 a_1522_3425.n1 a_1522_3425.n0 173.817
R18933 a_1522_3425.n1 a_1522_3425.t1 20.826
R18934 a_1522_3425.n2 a_1522_3425.n1 20.689
R18935 a_1892_3425.t0 a_1892_3425.t1 242.857
R18936 a_6697_975.n0 a_6697_975.t2 358.166
R18937 a_6697_975.t5 a_6697_975.t3 337.399
R18938 a_6697_975.t3 a_6697_975.t4 285.986
R18939 a_6697_975.n0 a_6697_975.t5 282.573
R18940 a_6697_975.n1 a_6697_975.t0 202.857
R18941 a_6697_975.n1 a_6697_975.n0 173.817
R18942 a_6697_975.n1 a_6697_975.t1 20.826
R18943 a_6697_975.n2 a_6697_975.n1 20.689
R18944 a_13934_n5338.n0 a_13934_n5338.t0 63.08
R18945 a_13934_n5338.n0 a_13934_n5338.t2 41.307
R18946 a_13934_n5338.t1 a_13934_n5338.n0 2.251
R18947 a_947_2180.n0 a_947_2180.t0 358.166
R18948 a_947_2180.t4 a_947_2180.t5 337.399
R18949 a_947_2180.t5 a_947_2180.t3 285.986
R18950 a_947_2180.n0 a_947_2180.t4 282.573
R18951 a_947_2180.n1 a_947_2180.t2 202.857
R18952 a_947_2180.n1 a_947_2180.n0 173.817
R18953 a_947_2180.n1 a_947_2180.t1 20.826
R18954 a_947_2180.n2 a_947_2180.n1 20.689
R18955 a_2672_1698.n0 a_2672_1698.t1 358.166
R18956 a_2672_1698.t3 a_2672_1698.t4 337.399
R18957 a_2672_1698.t4 a_2672_1698.t5 285.986
R18958 a_2672_1698.n0 a_2672_1698.t3 282.573
R18959 a_2672_1698.n1 a_2672_1698.t0 202.857
R18960 a_2672_1698.n1 a_2672_1698.n0 173.817
R18961 a_2672_1698.n1 a_2672_1698.t2 20.826
R18962 a_2672_1698.n2 a_2672_1698.n1 20.689
R18963 a_2577_1683.n0 a_2577_1683.t1 362.857
R18964 a_2577_1683.t3 a_2577_1683.t4 337.399
R18965 a_2577_1683.t4 a_2577_1683.t5 298.839
R18966 a_2577_1683.n0 a_2577_1683.t3 280.405
R18967 a_2577_1683.n1 a_2577_1683.t2 200
R18968 a_2577_1683.n1 a_2577_1683.n0 172.311
R18969 a_2577_1683.n2 a_2577_1683.n1 24
R18970 a_2577_1683.n1 a_2577_1683.t0 21.212
R18971 a_7752_n1068.n0 a_7752_n1068.t2 362.857
R18972 a_7752_n1068.t4 a_7752_n1068.t5 337.399
R18973 a_7752_n1068.t5 a_7752_n1068.t3 298.839
R18974 a_7752_n1068.n0 a_7752_n1068.t4 280.405
R18975 a_7752_n1068.n1 a_7752_n1068.t0 200
R18976 a_7752_n1068.n1 a_7752_n1068.n0 172.311
R18977 a_7752_n1068.n2 a_7752_n1068.n1 24
R18978 a_7752_n1068.n1 a_7752_n1068.t1 21.212
R18979 a_4315_2180.t0 a_4315_2180.t1 242.857
R18980 a_7190_1216.t0 a_7190_1216.t1 242.857
R18981 a_6027_196.n0 a_6027_196.t1 362.857
R18982 a_6027_196.t4 a_6027_196.t3 337.399
R18983 a_6027_196.t3 a_6027_196.t5 298.839
R18984 a_6027_196.n0 a_6027_196.t4 280.405
R18985 a_6027_196.n1 a_6027_196.t2 200
R18986 a_6027_196.n1 a_6027_196.n0 172.311
R18987 a_6027_196.n2 a_6027_196.n1 24
R18988 a_6027_196.n1 a_6027_196.t0 21.212
R18989 a_5547_3666.n0 a_5547_3666.t1 358.166
R18990 a_5547_3666.t4 a_5547_3666.t5 337.399
R18991 a_5547_3666.t5 a_5547_3666.t3 285.986
R18992 a_5547_3666.n0 a_5547_3666.t4 282.573
R18993 a_5547_3666.n1 a_5547_3666.t2 202.857
R18994 a_5547_3666.n1 a_5547_3666.n0 173.817
R18995 a_5547_3666.n1 a_5547_3666.t0 20.826
R18996 a_5547_3666.n2 a_5547_3666.n1 20.689
R18997 a_5917_3666.t0 a_5917_3666.t1 242.857
R18998 a_7752_678.n0 a_7752_678.t2 362.857
R18999 a_7752_678.t4 a_7752_678.t3 337.399
R19000 a_7752_678.t3 a_7752_678.t5 298.839
R19001 a_7752_678.n0 a_7752_678.t4 280.405
R19002 a_7752_678.n1 a_7752_678.t0 200
R19003 a_7752_678.n1 a_7752_678.n0 172.311
R19004 a_7752_678.n2 a_7752_678.n1 24
R19005 a_7752_678.n1 a_7752_678.t1 21.212
R19006 a_7847_693.n0 a_7847_693.t1 358.166
R19007 a_7847_693.t5 a_7847_693.t4 337.399
R19008 a_7847_693.t4 a_7847_693.t3 285.986
R19009 a_7847_693.n0 a_7847_693.t5 282.573
R19010 a_7847_693.n1 a_7847_693.t2 202.857
R19011 a_7847_693.n1 a_7847_693.n0 173.817
R19012 a_7847_693.n1 a_7847_693.t0 20.826
R19013 a_7847_693.n2 a_7847_693.n1 20.689
R19014 a_4745_n5338.n0 a_4745_n5338.t0 63.08
R19015 a_4745_n5338.n0 a_4745_n5338.t2 41.307
R19016 a_4745_n5338.t1 a_4745_n5338.n0 2.251
R19017 a_4883_n5338.t0 a_4883_n5338.t1 68.74
R19018 a_2672_n812.n0 a_2672_n812.t2 358.166
R19019 a_2672_n812.t3 a_2672_n812.t4 337.399
R19020 a_2672_n812.t4 a_2672_n812.t5 285.986
R19021 a_2672_n812.n0 a_2672_n812.t3 282.573
R19022 a_2672_n812.n1 a_2672_n812.t0 202.857
R19023 a_2672_n812.n1 a_2672_n812.n0 173.817
R19024 a_2672_n812.n1 a_2672_n812.t1 20.826
R19025 a_2672_n812.n2 a_2672_n812.n1 20.689
R19026 a_2577_n827.n0 a_2577_n827.t2 362.857
R19027 a_2577_n827.t5 a_2577_n827.t3 337.399
R19028 a_2577_n827.t3 a_2577_n827.t4 298.839
R19029 a_2577_n827.n0 a_2577_n827.t5 280.405
R19030 a_2577_n827.n1 a_2577_n827.t0 200
R19031 a_2577_n827.n1 a_2577_n827.n0 172.311
R19032 a_2577_n827.n2 a_2577_n827.n1 24
R19033 a_2577_n827.n1 a_2577_n827.t1 21.212
R19034 a_4302_4133.n0 a_4302_4133.t2 362.857
R19035 a_4302_4133.t3 a_4302_4133.t5 337.399
R19036 a_4302_4133.t5 a_4302_4133.t4 298.839
R19037 a_4302_4133.n0 a_4302_4133.t3 280.405
R19038 a_4302_4133.n1 a_4302_4133.t1 200
R19039 a_4302_4133.n1 a_4302_4133.n0 172.311
R19040 a_4302_4133.n2 a_4302_4133.n1 24
R19041 a_4302_4133.n1 a_4302_4133.t0 21.212
R19042 a_4397_4148.n0 a_4397_4148.t2 358.166
R19043 a_4397_4148.t5 a_4397_4148.t3 337.399
R19044 a_4397_4148.t3 a_4397_4148.t4 285.986
R19045 a_4397_4148.n0 a_4397_4148.t5 282.573
R19046 a_4397_4148.n1 a_4397_4148.t0 202.857
R19047 a_4397_4148.n1 a_4397_4148.n0 173.817
R19048 a_4397_4148.n1 a_4397_4148.t1 20.826
R19049 a_4397_4148.n2 a_4397_4148.n1 20.689
R19050 a_5452_2165.n0 a_5452_2165.t1 362.857
R19051 a_5452_2165.t3 a_5452_2165.t4 337.399
R19052 a_5452_2165.t4 a_5452_2165.t5 298.839
R19053 a_5452_2165.n0 a_5452_2165.t3 280.405
R19054 a_5452_2165.n1 a_5452_2165.t0 200
R19055 a_5452_2165.n1 a_5452_2165.n0 172.311
R19056 a_5452_2165.n2 a_5452_2165.n1 24
R19057 a_5452_2165.n1 a_5452_2165.t2 21.212
R19058 a_5547_2180.n0 a_5547_2180.t2 358.166
R19059 a_5547_2180.t4 a_5547_2180.t5 337.399
R19060 a_5547_2180.t5 a_5547_2180.t3 285.986
R19061 a_5547_2180.n0 a_5547_2180.t4 282.573
R19062 a_5547_2180.n1 a_5547_2180.t0 202.857
R19063 a_5547_2180.n1 a_5547_2180.n0 173.817
R19064 a_5547_2180.n1 a_5547_2180.t1 20.826
R19065 a_5547_2180.n2 a_5547_2180.n1 20.689
R19066 a_3995_4887.n25 a_3995_4887.t27 561.971
R19067 a_3995_4887.n0 a_3995_4887.t6 449.944
R19068 a_3995_4887.t15 a_3995_4887.n25 108.636
R19069 a_3995_4887.n0 a_3995_4887.t5 74.821
R19070 a_3995_4887.n24 a_3995_4887.t22 63.519
R19071 a_3995_4887.n23 a_3995_4887.t1 63.519
R19072 a_3995_4887.n22 a_3995_4887.t14 63.519
R19073 a_3995_4887.n21 a_3995_4887.t16 63.519
R19074 a_3995_4887.n20 a_3995_4887.t13 63.519
R19075 a_3995_4887.n19 a_3995_4887.t19 63.519
R19076 a_3995_4887.n18 a_3995_4887.t20 63.519
R19077 a_3995_4887.n17 a_3995_4887.t10 63.519
R19078 a_3995_4887.n16 a_3995_4887.t4 63.519
R19079 a_3995_4887.n15 a_3995_4887.t8 63.519
R19080 a_3995_4887.n14 a_3995_4887.t23 63.519
R19081 a_3995_4887.n13 a_3995_4887.t21 63.519
R19082 a_3995_4887.n12 a_3995_4887.t18 63.519
R19083 a_3995_4887.n11 a_3995_4887.t11 63.519
R19084 a_3995_4887.n10 a_3995_4887.t12 63.519
R19085 a_3995_4887.n9 a_3995_4887.t24 63.519
R19086 a_3995_4887.n8 a_3995_4887.t0 63.519
R19087 a_3995_4887.n7 a_3995_4887.t3 63.519
R19088 a_3995_4887.n6 a_3995_4887.t2 63.519
R19089 a_3995_4887.n5 a_3995_4887.t26 63.519
R19090 a_3995_4887.n4 a_3995_4887.t9 63.519
R19091 a_3995_4887.n3 a_3995_4887.t17 63.519
R19092 a_3995_4887.n2 a_3995_4887.t25 63.519
R19093 a_3995_4887.n1 a_3995_4887.t7 63.519
R19094 a_3995_4887.n1 a_3995_4887.n0 8.619
R19095 a_3995_4887.n25 a_3995_4887.n24 2.946
R19096 a_3995_4887.n23 a_3995_4887.n22 2.524
R19097 a_3995_4887.n3 a_3995_4887.n2 2.498
R19098 a_3995_4887.n17 a_3995_4887.n16 2.364
R19099 a_3995_4887.n9 a_3995_4887.n8 2.355
R19100 a_3995_4887.n24 a_3995_4887.n23 1.998
R19101 a_3995_4887.n22 a_3995_4887.n21 1.998
R19102 a_3995_4887.n21 a_3995_4887.n20 1.998
R19103 a_3995_4887.n20 a_3995_4887.n19 1.998
R19104 a_3995_4887.n19 a_3995_4887.n18 1.998
R19105 a_3995_4887.n18 a_3995_4887.n17 1.998
R19106 a_3995_4887.n16 a_3995_4887.n15 1.998
R19107 a_3995_4887.n15 a_3995_4887.n14 1.998
R19108 a_3995_4887.n14 a_3995_4887.n13 1.998
R19109 a_3995_4887.n13 a_3995_4887.n12 1.998
R19110 a_3995_4887.n12 a_3995_4887.n11 1.998
R19111 a_3995_4887.n11 a_3995_4887.n10 1.998
R19112 a_3995_4887.n10 a_3995_4887.n9 1.998
R19113 a_3995_4887.n8 a_3995_4887.n7 1.998
R19114 a_3995_4887.n7 a_3995_4887.n6 1.998
R19115 a_3995_4887.n6 a_3995_4887.n5 1.998
R19116 a_3995_4887.n5 a_3995_4887.n4 1.998
R19117 a_3995_4887.n4 a_3995_4887.n3 1.998
R19118 a_3995_4887.n2 a_3995_4887.n1 1.998
R19119 a_3727_1442.n0 a_3727_1442.t1 362.857
R19120 a_3727_1442.t5 a_3727_1442.t3 337.399
R19121 a_3727_1442.t3 a_3727_1442.t4 298.839
R19122 a_3727_1442.n0 a_3727_1442.t5 280.405
R19123 a_3727_1442.n1 a_3727_1442.t2 200
R19124 a_3727_1442.n1 a_3727_1442.n0 172.311
R19125 a_3727_1442.n2 a_3727_1442.n1 24
R19126 a_3727_1442.n1 a_3727_1442.t0 21.212
R19127 a_5547_n512.n0 a_5547_n512.t1 358.166
R19128 a_5547_n512.t5 a_5547_n512.t3 337.399
R19129 a_5547_n512.t3 a_5547_n512.t4 285.986
R19130 a_5547_n512.n0 a_5547_n512.t5 282.573
R19131 a_5547_n512.n1 a_5547_n512.t0 202.857
R19132 a_5547_n512.n1 a_5547_n512.n0 173.817
R19133 a_5547_n512.n1 a_5547_n512.t2 20.826
R19134 a_5547_n512.n2 a_5547_n512.n1 20.689
R19135 a_5452_n527.n0 a_5452_n527.t1 362.857
R19136 a_5452_n527.t3 a_5452_n527.t4 337.399
R19137 a_5452_n527.t4 a_5452_n527.t5 298.839
R19138 a_5452_n527.n0 a_5452_n527.t3 280.405
R19139 a_5452_n527.n1 a_5452_n527.t2 200
R19140 a_5452_n527.n1 a_5452_n527.n0 172.311
R19141 a_5452_n527.n2 a_5452_n527.n1 24
R19142 a_5452_n527.n1 a_5452_n527.t0 21.212
R19143 a_865_452.t0 a_865_452.t1 242.857
R19144 a_7272_1698.n0 a_7272_1698.t0 358.166
R19145 a_7272_1698.t4 a_7272_1698.t3 337.399
R19146 a_7272_1698.t3 a_7272_1698.t5 285.986
R19147 a_7272_1698.n0 a_7272_1698.t4 282.573
R19148 a_7272_1698.n1 a_7272_1698.t1 202.857
R19149 a_7272_1698.n1 a_7272_1698.n0 173.817
R19150 a_7272_1698.n1 a_7272_1698.t2 20.826
R19151 a_7272_1698.n2 a_7272_1698.n1 20.689
R19152 a_7177_1683.n0 a_7177_1683.t2 362.857
R19153 a_7177_1683.t5 a_7177_1683.t3 337.399
R19154 a_7177_1683.t3 a_7177_1683.t4 298.839
R19155 a_7177_1683.n0 a_7177_1683.t5 280.405
R19156 a_7177_1683.n1 a_7177_1683.t0 200
R19157 a_7177_1683.n1 a_7177_1683.n0 172.311
R19158 a_7177_1683.n2 a_7177_1683.n1 24
R19159 a_7177_1683.n1 a_7177_1683.t1 21.212
R19160 a_6268_n2426.n3 a_6268_n2426.t3 475.39
R19161 a_6268_n2426.n3 a_6268_n2426.n2 365.296
R19162 a_6268_n2426.t5 a_6268_n2426.t7 228.696
R19163 a_6268_n2426.n2 a_6268_n2426.t1 185.704
R19164 a_6268_n2426.n0 a_6268_n2426.t5 126.761
R19165 a_6268_n2426.n1 a_6268_n2426.t6 126.284
R19166 a_6268_n2426.n1 a_6268_n2426.t0 126.284
R19167 a_6268_n2426.t2 a_6268_n2426.n3 124.375
R19168 a_6268_n2426.t0 a_6268_n2426.n0 115.122
R19169 a_6268_n2426.n0 a_6268_n2426.t4 111.229
R19170 a_6268_n2426.n2 a_6268_n2426.n1 8.764
R19171 a_7959_n5092.t0 a_7959_n5092.t1 42.705
R19172 a_7109_n5338.n0 a_7109_n5338.t0 63.08
R19173 a_7109_n5338.n0 a_7109_n5338.t2 41.307
R19174 a_7109_n5338.t1 a_7109_n5338.n0 2.251
R19175 a_7247_n5338.t0 a_7247_n5338.t1 68.74
R19176 a_3822_1216.n0 a_3822_1216.t1 358.166
R19177 a_3822_1216.t4 a_3822_1216.t3 337.399
R19178 a_3822_1216.t3 a_3822_1216.t5 285.986
R19179 a_3822_1216.n0 a_3822_1216.t4 282.573
R19180 a_3822_1216.n1 a_3822_1216.t0 202.857
R19181 a_3822_1216.n1 a_3822_1216.n0 173.817
R19182 a_3822_1216.n1 a_3822_1216.t2 20.826
R19183 a_3822_1216.n2 a_3822_1216.n1 20.689
R19184 a_3727_1201.n0 a_3727_1201.t1 362.857
R19185 a_3727_1201.t3 a_3727_1201.t4 337.399
R19186 a_3727_1201.t4 a_3727_1201.t5 298.839
R19187 a_3727_1201.n0 a_3727_1201.t3 280.405
R19188 a_3727_1201.n1 a_3727_1201.t2 200
R19189 a_3727_1201.n1 a_3727_1201.n0 172.311
R19190 a_3727_1201.n2 a_3727_1201.n1 24
R19191 a_3727_1201.n1 a_3727_1201.t0 21.212
R19192 a_3617_975.t0 a_3617_975.t1 242.857
R19193 a_7418_n2426.n3 a_7418_n2426.t3 475.39
R19194 a_7418_n2426.n3 a_7418_n2426.n2 273.59
R19195 a_7418_n2426.t5 a_7418_n2426.t7 228.696
R19196 a_7418_n2426.n2 a_7418_n2426.t1 185.704
R19197 a_7418_n2426.n0 a_7418_n2426.t5 126.761
R19198 a_7418_n2426.n1 a_7418_n2426.t6 126.284
R19199 a_7418_n2426.n1 a_7418_n2426.t0 126.284
R19200 a_7418_n2426.t2 a_7418_n2426.n3 124.375
R19201 a_7418_n2426.t0 a_7418_n2426.n0 115.122
R19202 a_7418_n2426.n0 a_7418_n2426.t4 111.229
R19203 a_7418_n2426.n2 a_7418_n2426.n1 8.764
R19204 a_10327_n5092.t0 a_10327_n5092.t1 42.705
R19205 a_9367_452.t0 a_9367_452.t1 242.857
R19206 a_7272_n812.n0 a_7272_n812.t1 358.166
R19207 a_7272_n812.t4 a_7272_n812.t3 337.399
R19208 a_7272_n812.t3 a_7272_n812.t5 285.986
R19209 a_7272_n812.n0 a_7272_n812.t4 282.573
R19210 a_7272_n812.n1 a_7272_n812.t0 202.857
R19211 a_7272_n812.n1 a_7272_n812.n0 173.817
R19212 a_7272_n812.n1 a_7272_n812.t2 20.826
R19213 a_7272_n812.n2 a_7272_n812.n1 20.689
R19214 a_7177_n827.n0 a_7177_n827.t2 362.857
R19215 a_7177_n827.t3 a_7177_n827.t4 337.399
R19216 a_7177_n827.t4 a_7177_n827.t5 298.839
R19217 a_7177_n827.n0 a_7177_n827.t3 280.405
R19218 a_7177_n827.n1 a_7177_n827.t0 200
R19219 a_7177_n827.n1 a_7177_n827.n0 172.311
R19220 a_7177_n827.n2 a_7177_n827.n1 24
R19221 a_7177_n827.n1 a_7177_n827.t1 21.212
R19222 a_5342_4445.t0 a_5342_4445.t1 242.857
R19223 a_7067_3907.t0 a_7067_3907.t1 242.857
R19224 a_1427_2647.n0 a_1427_2647.t1 362.857
R19225 a_1427_2647.t5 a_1427_2647.t3 337.399
R19226 a_1427_2647.t3 a_1427_2647.t4 298.839
R19227 a_1427_2647.n0 a_1427_2647.t5 280.405
R19228 a_1427_2647.n1 a_1427_2647.t2 200
R19229 a_1427_2647.n1 a_1427_2647.n0 172.311
R19230 a_1427_2647.n2 a_1427_2647.n1 24
R19231 a_1427_2647.n1 a_1427_2647.t0 21.212
R19232 a_1522_2662.n0 a_1522_2662.t1 358.166
R19233 a_1522_2662.t4 a_1522_2662.t3 337.399
R19234 a_1522_2662.t3 a_1522_2662.t5 285.986
R19235 a_1522_2662.n0 a_1522_2662.t4 282.573
R19236 a_1522_2662.n1 a_1522_2662.t2 202.857
R19237 a_1522_2662.n1 a_1522_2662.n0 173.817
R19238 a_1522_2662.n1 a_1522_2662.t0 20.826
R19239 a_1522_2662.n2 a_1522_2662.n1 20.689
R19240 a_2097_2180.n0 a_2097_2180.t2 358.166
R19241 a_2097_2180.t4 a_2097_2180.t5 337.399
R19242 a_2097_2180.t5 a_2097_2180.t3 285.986
R19243 a_2097_2180.n0 a_2097_2180.t4 282.573
R19244 a_2097_2180.n1 a_2097_2180.t0 202.857
R19245 a_2097_2180.n1 a_2097_2180.n0 173.817
R19246 a_2097_2180.n1 a_2097_2180.t1 20.826
R19247 a_2097_2180.n2 a_2097_2180.n1 20.689
R19248 a_8327_678.n0 a_8327_678.t2 362.857
R19249 a_8327_678.t5 a_8327_678.t4 337.399
R19250 a_8327_678.t4 a_8327_678.t3 298.839
R19251 a_8327_678.n0 a_8327_678.t5 280.405
R19252 a_8327_678.n1 a_8327_678.t1 200
R19253 a_8327_678.n1 a_8327_678.n0 172.311
R19254 a_8327_678.n2 a_8327_678.n1 24
R19255 a_8327_678.n1 a_8327_678.t0 21.212
R19256 a_8340_693.t0 a_8340_693.t1 242.857
R19257 a_5452_n45.n0 a_5452_n45.t1 362.857
R19258 a_5452_n45.t3 a_5452_n45.t5 337.399
R19259 a_5452_n45.t5 a_5452_n45.t4 298.839
R19260 a_5452_n45.n0 a_5452_n45.t3 280.405
R19261 a_5452_n45.n1 a_5452_n45.t0 200
R19262 a_5452_n45.n1 a_5452_n45.n0 172.311
R19263 a_5452_n45.n2 a_5452_n45.n1 24
R19264 a_5452_n45.n1 a_5452_n45.t2 21.212
R19265 a_5547_n30.n0 a_5547_n30.t2 358.166
R19266 a_5547_n30.t3 a_5547_n30.t5 337.399
R19267 a_5547_n30.t5 a_5547_n30.t4 285.986
R19268 a_5547_n30.n0 a_5547_n30.t3 282.573
R19269 a_5547_n30.n1 a_5547_n30.t0 202.857
R19270 a_5547_n30.n1 a_5547_n30.n0 173.817
R19271 a_5547_n30.n1 a_5547_n30.t1 20.826
R19272 a_5547_n30.n2 a_5547_n30.n1 20.689
R19273 a_2672_4686.n0 a_2672_4686.t1 358.166
R19274 a_2672_4686.t5 a_2672_4686.t3 337.399
R19275 a_2672_4686.t3 a_2672_4686.t4 285.986
R19276 a_2672_4686.n0 a_2672_4686.t5 282.573
R19277 a_2672_4686.n1 a_2672_4686.t0 202.857
R19278 a_2672_4686.n1 a_2672_4686.n0 173.817
R19279 a_2672_4686.n1 a_2672_4686.t2 20.826
R19280 a_2672_4686.n2 a_2672_4686.n1 20.689
R19281 a_2577_4671.n0 a_2577_4671.t2 362.857
R19282 a_2577_4671.t5 a_2577_4671.t3 337.399
R19283 a_2577_4671.t3 a_2577_4671.t4 298.839
R19284 a_2577_4671.n0 a_2577_4671.t5 280.405
R19285 a_2577_4671.n1 a_2577_4671.t0 200
R19286 a_2577_4671.n1 a_2577_4671.n0 172.311
R19287 a_2577_4671.n2 a_2577_4671.n1 24
R19288 a_2577_4671.n1 a_2577_4671.t1 21.212
R19289 a_6615_4445.t0 a_6615_4445.t1 242.857
R19290 a_5630_n3770.n0 a_5630_n3770.t0 65.064
R19291 a_5630_n3770.n0 a_5630_n3770.t2 42.011
R19292 a_5630_n3770.t1 a_5630_n3770.n0 2.113
R19293 a_6602_1201.n0 a_6602_1201.t1 362.857
R19294 a_6602_1201.t3 a_6602_1201.t5 337.399
R19295 a_6602_1201.t5 a_6602_1201.t4 298.839
R19296 a_6602_1201.n0 a_6602_1201.t3 280.405
R19297 a_6602_1201.n1 a_6602_1201.t2 200
R19298 a_6602_1201.n1 a_6602_1201.n0 172.311
R19299 a_6602_1201.n2 a_6602_1201.n1 24
R19300 a_6602_1201.n1 a_6602_1201.t0 21.212
R19301 a_1522_n512.n0 a_1522_n512.t1 358.166
R19302 a_1522_n512.t3 a_1522_n512.t5 337.399
R19303 a_1522_n512.t5 a_1522_n512.t4 285.986
R19304 a_1522_n512.n0 a_1522_n512.t3 282.573
R19305 a_1522_n512.n1 a_1522_n512.t2 202.857
R19306 a_1522_n512.n1 a_1522_n512.n0 173.817
R19307 a_1522_n512.n1 a_1522_n512.t0 20.826
R19308 a_1522_n512.n2 a_1522_n512.n1 20.689
R19309 a_3328_n2086.t0 a_3328_n2086.t1 34.8
R19310 a_852_n1068.n0 a_852_n1068.t1 362.857
R19311 a_852_n1068.t5 a_852_n1068.t3 337.399
R19312 a_852_n1068.t3 a_852_n1068.t4 298.839
R19313 a_852_n1068.n0 a_852_n1068.t5 280.405
R19314 a_852_n1068.n1 a_852_n1068.t0 200
R19315 a_852_n1068.n1 a_852_n1068.n0 172.311
R19316 a_852_n1068.n2 a_852_n1068.n1 24
R19317 a_852_n1068.n1 a_852_n1068.t2 21.212
R19318 a_947_n1053.n0 a_947_n1053.t1 358.166
R19319 a_947_n1053.t4 a_947_n1053.t5 337.399
R19320 a_947_n1053.t5 a_947_n1053.t3 285.986
R19321 a_947_n1053.n0 a_947_n1053.t4 282.573
R19322 a_947_n1053.n1 a_947_n1053.t2 202.857
R19323 a_947_n1053.n1 a_947_n1053.n0 173.817
R19324 a_947_n1053.n1 a_947_n1053.t0 20.826
R19325 a_947_n1053.n2 a_947_n1053.n1 20.689
R19326 a_372_4148.n0 a_372_4148.t0 358.166
R19327 a_372_4148.t3 a_372_4148.t5 337.399
R19328 a_372_4148.t5 a_372_4148.t4 285.986
R19329 a_372_4148.n0 a_372_4148.t3 282.573
R19330 a_372_4148.n1 a_372_4148.t2 202.857
R19331 a_372_4148.n1 a_372_4148.n0 173.817
R19332 a_372_4148.n1 a_372_4148.t1 20.826
R19333 a_372_4148.n2 a_372_4148.n1 20.689
R19334 a_7752_2647.n0 a_7752_2647.t2 362.857
R19335 a_7752_2647.t4 a_7752_2647.t5 337.399
R19336 a_7752_2647.t5 a_7752_2647.t3 298.839
R19337 a_7752_2647.n0 a_7752_2647.t4 280.405
R19338 a_7752_2647.n1 a_7752_2647.t0 200
R19339 a_7752_2647.n1 a_7752_2647.n0 172.311
R19340 a_7752_2647.n2 a_7752_2647.n1 24
R19341 a_7752_2647.n1 a_7752_2647.t1 21.212
R19342 a_7765_2662.t0 a_7765_2662.t1 242.857
R19343 a_2672_1216.n0 a_2672_1216.t0 358.166
R19344 a_2672_1216.t3 a_2672_1216.t4 337.399
R19345 a_2672_1216.t4 a_2672_1216.t5 285.986
R19346 a_2672_1216.n0 a_2672_1216.t3 282.573
R19347 a_2672_1216.n1 a_2672_1216.t1 202.857
R19348 a_2672_1216.n1 a_2672_1216.n0 173.817
R19349 a_2672_1216.n1 a_2672_1216.t2 20.826
R19350 a_2672_1216.n2 a_2672_1216.n1 20.689
R19351 a_2577_1201.n0 a_2577_1201.t2 362.857
R19352 a_2577_1201.t3 a_2577_1201.t4 337.399
R19353 a_2577_1201.t4 a_2577_1201.t5 298.839
R19354 a_2577_1201.n0 a_2577_1201.t3 280.405
R19355 a_2577_1201.n1 a_2577_1201.t0 200
R19356 a_2577_1201.n1 a_2577_1201.n0 172.311
R19357 a_2577_1201.n2 a_2577_1201.n1 24
R19358 a_2577_1201.n1 a_2577_1201.t1 21.212
R19359 a_8221_n4483.n0 a_8221_n4483.t3 1464.36
R19360 a_8221_n4483.n0 a_8221_n4483.t4 713.588
R19361 a_8221_n4483.n1 a_8221_n4483.t0 374.998
R19362 a_8221_n4483.n1 a_8221_n4483.t2 273.351
R19363 a_8221_n4483.n2 a_8221_n4483.n0 143.764
R19364 a_8221_n4483.t1 a_8221_n4483.n2 78.209
R19365 a_8221_n4483.n2 a_8221_n4483.n1 4.517
R19366 ADC10_OUT[0].n0 ADC10_OUT[0].t3 1354.27
R19367 ADC10_OUT[0].n0 ADC10_OUT[0].t4 821.954
R19368 ADC10_OUT[0].n3 ADC10_OUT[0].t0 334.338
R19369 ADC10_OUT[0].n2 ADC10_OUT[0].t1 266.575
R19370 ADC10_OUT[0].n1 ADC10_OUT[0].n0 149.035
R19371 ADC10_OUT[0] ADC10_OUT[0].n3 61.901
R19372 ADC10_OUT[0].n3 ADC10_OUT[0].n2 49.694
R19373 ADC10_OUT[0].n1 ADC10_OUT[0].t2 46.723
R19374 ADC10_OUT[0].n2 ADC10_OUT[0].n1 17.317
R19375 a_7994_n3770.n0 a_7994_n3770.t0 65.064
R19376 a_7994_n3770.n0 a_7994_n3770.t2 42.011
R19377 a_7994_n3770.t1 a_7994_n3770.n0 2.113
R19378 a_10589_n7216.n0 a_10589_n7216.t3 1464.36
R19379 a_10589_n7216.n0 a_10589_n7216.t4 713.588
R19380 a_10589_n7216.n1 a_10589_n7216.t0 374.998
R19381 a_10589_n7216.n1 a_10589_n7216.t2 273.351
R19382 a_10589_n7216.n2 a_10589_n7216.n0 143.764
R19383 a_10589_n7216.t1 a_10589_n7216.n2 78.209
R19384 a_10589_n7216.n2 a_10589_n7216.n1 4.517
R19385 a_10362_n6503.n0 a_10362_n6503.t1 65.064
R19386 a_10362_n6503.t0 a_10362_n6503.n0 42.011
R19387 a_10362_n6503.n0 a_10362_n6503.t2 2.113
R19388 a_3247_4445.n0 a_3247_4445.t1 358.166
R19389 a_3247_4445.t5 a_3247_4445.t3 337.399
R19390 a_3247_4445.t3 a_3247_4445.t4 285.986
R19391 a_3247_4445.n0 a_3247_4445.t5 282.573
R19392 a_3247_4445.n1 a_3247_4445.t0 202.857
R19393 a_3247_4445.n1 a_3247_4445.n0 173.817
R19394 a_3247_4445.n1 a_3247_4445.t2 20.826
R19395 a_3247_4445.n2 a_3247_4445.n1 20.689
R19396 a_3152_4430.n0 a_3152_4430.t1 362.857
R19397 a_3152_4430.t3 a_3152_4430.t4 337.399
R19398 a_3152_4430.t4 a_3152_4430.t5 298.839
R19399 a_3152_4430.n0 a_3152_4430.t3 280.405
R19400 a_3152_4430.n1 a_3152_4430.t2 200
R19401 a_3152_4430.n1 a_3152_4430.n0 172.311
R19402 a_3152_4430.n2 a_3152_4430.n1 24
R19403 a_3152_4430.n1 a_3152_4430.t0 21.212
R19404 a_6677_n2234.n2 a_6677_n2234.t1 282.97
R19405 a_6677_n2234.n1 a_6677_n2234.t4 240.683
R19406 a_6677_n2234.n0 a_6677_n2234.t2 209.208
R19407 a_6677_n2234.n0 a_6677_n2234.t3 194.167
R19408 a_6677_n2234.t0 a_6677_n2234.n2 183.404
R19409 a_6677_n2234.n1 a_6677_n2234.n0 14.805
R19410 a_6677_n2234.n2 a_6677_n2234.n1 6.415
R19411 a_6800_n2132.n0 a_6800_n2132.t2 489.336
R19412 a_6800_n2132.n0 a_6800_n2132.t1 243.258
R19413 a_6800_n2132.t0 a_6800_n2132.n0 214.415
R19414 a_6122_3666.n0 a_6122_3666.t1 358.166
R19415 a_6122_3666.t5 a_6122_3666.t4 337.399
R19416 a_6122_3666.t4 a_6122_3666.t3 285.986
R19417 a_6122_3666.n0 a_6122_3666.t5 282.573
R19418 a_6122_3666.n1 a_6122_3666.t2 202.857
R19419 a_6122_3666.n1 a_6122_3666.n0 173.817
R19420 a_6122_3666.n1 a_6122_3666.t0 20.826
R19421 a_6122_3666.n2 a_6122_3666.n1 20.689
R19422 a_6492_3666.t0 a_6492_3666.t1 242.857
R19423 a_7177_1924.n0 a_7177_1924.t2 362.857
R19424 a_7177_1924.t3 a_7177_1924.t4 337.399
R19425 a_7177_1924.t4 a_7177_1924.t5 298.839
R19426 a_7177_1924.n0 a_7177_1924.t3 280.405
R19427 a_7177_1924.n1 a_7177_1924.t0 200
R19428 a_7177_1924.n1 a_7177_1924.n0 172.311
R19429 a_7177_1924.n2 a_7177_1924.n1 24
R19430 a_7177_1924.n1 a_7177_1924.t1 21.212
R19431 a_6122_n512.n0 a_6122_n512.t2 358.166
R19432 a_6122_n512.t4 a_6122_n512.t3 337.399
R19433 a_6122_n512.t3 a_6122_n512.t5 285.986
R19434 a_6122_n512.n0 a_6122_n512.t4 282.573
R19435 a_6122_n512.n1 a_6122_n512.t0 202.857
R19436 a_6122_n512.n1 a_6122_n512.n0 173.817
R19437 a_6122_n512.n1 a_6122_n512.t1 20.826
R19438 a_6122_n512.n2 a_6122_n512.n1 20.689
R19439 a_6027_n527.n0 a_6027_n527.t1 362.857
R19440 a_6027_n527.t3 a_6027_n527.t4 337.399
R19441 a_6027_n527.t4 a_6027_n527.t5 298.839
R19442 a_6027_n527.n0 a_6027_n527.t3 280.405
R19443 a_6027_n527.n1 a_6027_n527.t2 200
R19444 a_6027_n527.n1 a_6027_n527.n0 172.311
R19445 a_6027_n527.n2 a_6027_n527.n1 24
R19446 a_6027_n527.n1 a_6027_n527.t0 21.212
R19447 a_3740_n512.t0 a_3740_n512.t1 242.857
R19448 RWL[13].n0 RWL[13].t1 154.243
R19449 RWL[13].n14 RWL[13].t14 149.249
R19450 RWL[13].n13 RWL[13].t11 149.249
R19451 RWL[13].n12 RWL[13].t9 149.249
R19452 RWL[13].n11 RWL[13].t3 149.249
R19453 RWL[13].n10 RWL[13].t13 149.249
R19454 RWL[13].n9 RWL[13].t5 149.249
R19455 RWL[13].n8 RWL[13].t4 149.249
R19456 RWL[13].n7 RWL[13].t15 149.249
R19457 RWL[13].n6 RWL[13].t6 149.249
R19458 RWL[13].n5 RWL[13].t0 149.249
R19459 RWL[13].n4 RWL[13].t8 149.249
R19460 RWL[13].n3 RWL[13].t7 149.249
R19461 RWL[13].n2 RWL[13].t12 149.249
R19462 RWL[13].n1 RWL[13].t10 149.249
R19463 RWL[13].n0 RWL[13].t2 149.249
R19464 RWL[13] RWL[13].n14 42.872
R19465 RWL[13].n1 RWL[13].n0 4.994
R19466 RWL[13].n2 RWL[13].n1 4.994
R19467 RWL[13].n3 RWL[13].n2 4.994
R19468 RWL[13].n4 RWL[13].n3 4.994
R19469 RWL[13].n5 RWL[13].n4 4.994
R19470 RWL[13].n6 RWL[13].n5 4.994
R19471 RWL[13].n7 RWL[13].n6 4.994
R19472 RWL[13].n8 RWL[13].n7 4.994
R19473 RWL[13].n9 RWL[13].n8 4.994
R19474 RWL[13].n10 RWL[13].n9 4.994
R19475 RWL[13].n11 RWL[13].n10 4.994
R19476 RWL[13].n12 RWL[13].n11 4.994
R19477 RWL[13].n13 RWL[13].n12 4.994
R19478 RWL[13].n14 RWL[13].n13 4.994
R19479 a_5465_452.t0 a_5465_452.t1 242.857
R19480 a_3042_3184.t0 a_3042_3184.t1 242.857
R19481 a_7272_1216.n0 a_7272_1216.t0 358.166
R19482 a_7272_1216.t4 a_7272_1216.t3 337.399
R19483 a_7272_1216.t3 a_7272_1216.t5 285.986
R19484 a_7272_1216.n0 a_7272_1216.t4 282.573
R19485 a_7272_1216.n1 a_7272_1216.t1 202.857
R19486 a_7272_1216.n1 a_7272_1216.n0 173.817
R19487 a_7272_1216.n1 a_7272_1216.t2 20.826
R19488 a_7272_1216.n2 a_7272_1216.n1 20.689
R19489 a_7177_1201.n0 a_7177_1201.t2 362.857
R19490 a_7177_1201.t5 a_7177_1201.t3 337.399
R19491 a_7177_1201.t3 a_7177_1201.t4 298.839
R19492 a_7177_1201.n0 a_7177_1201.t5 280.405
R19493 a_7177_1201.n1 a_7177_1201.t0 200
R19494 a_7177_1201.n1 a_7177_1201.n0 172.311
R19495 a_7177_1201.n2 a_7177_1201.n1 24
R19496 a_7177_1201.n1 a_7177_1201.t1 21.212
R19497 a_8217_693.t0 a_8217_693.t1 242.857
R19498 ADC12_OUT[0].n0 ADC12_OUT[0].t4 1354.27
R19499 ADC12_OUT[0].n0 ADC12_OUT[0].t3 821.954
R19500 ADC12_OUT[0].n3 ADC12_OUT[0].t0 339.609
R19501 ADC12_OUT[0].n2 ADC12_OUT[0].t2 266.575
R19502 ADC12_OUT[0].n1 ADC12_OUT[0].n0 149.035
R19503 ADC12_OUT[0] ADC12_OUT[0].n3 61.776
R19504 ADC12_OUT[0].n1 ADC12_OUT[0].t1 46.723
R19505 ADC12_OUT[0].n3 ADC12_OUT[0].n2 44.423
R19506 ADC12_OUT[0].n2 ADC12_OUT[0].n1 17.317
R19507 a_10589_n4483.n0 a_10589_n4483.t3 1464.36
R19508 a_10589_n4483.n0 a_10589_n4483.t4 713.588
R19509 a_10589_n4483.n1 a_10589_n4483.t0 374.998
R19510 a_10589_n4483.n1 a_10589_n4483.t2 273.351
R19511 a_10589_n4483.n2 a_10589_n4483.n0 143.764
R19512 a_10589_n4483.t1 a_10589_n4483.n2 78.209
R19513 a_10589_n4483.n2 a_10589_n4483.n1 4.517
R19514 a_7067_n271.t0 a_7067_n271.t1 242.857
R19515 ADC1_OUT[3].n0 ADC1_OUT[3].t4 1355.37
R19516 ADC1_OUT[3].n0 ADC1_OUT[3].t3 820.859
R19517 ADC1_OUT[3].n3 ADC1_OUT[3].t0 331.396
R19518 ADC1_OUT[3].n2 ADC1_OUT[3].t1 266.644
R19519 ADC1_OUT[3].n1 ADC1_OUT[3].n0 149.035
R19520 ADC1_OUT[3].n3 ADC1_OUT[3].n2 52.705
R19521 ADC1_OUT[3].n1 ADC1_OUT[3].t2 45.968
R19522 ADC1_OUT[3] ADC1_OUT[3].n3 22.338
R19523 ADC1_OUT[3].n2 ADC1_OUT[3].n1 17.317
R19524 a_n2415_n8583.n0 a_n2415_n8583.t3 1465.51
R19525 a_n2415_n8583.n0 a_n2415_n8583.t4 712.44
R19526 a_n2415_n8583.n1 a_n2415_n8583.t0 375.067
R19527 a_n2415_n8583.n1 a_n2415_n8583.t1 272.668
R19528 a_n2415_n8583.n2 a_n2415_n8583.n0 143.764
R19529 a_n2415_n8583.t2 a_n2415_n8583.n2 78.193
R19530 a_n2415_n8583.n2 a_n2415_n8583.n1 4.517
R19531 a_7272_n1053.n0 a_7272_n1053.t2 358.166
R19532 a_7272_n1053.t3 a_7272_n1053.t5 337.399
R19533 a_7272_n1053.t5 a_7272_n1053.t4 285.986
R19534 a_7272_n1053.n0 a_7272_n1053.t3 282.573
R19535 a_7272_n1053.n1 a_7272_n1053.t0 202.857
R19536 a_7272_n1053.n1 a_7272_n1053.n0 173.817
R19537 a_7272_n1053.n1 a_7272_n1053.t1 20.826
R19538 a_7272_n1053.n2 a_7272_n1053.n1 20.689
R19539 a_7177_n1068.n0 a_7177_n1068.t2 362.857
R19540 a_7177_n1068.t5 a_7177_n1068.t3 337.399
R19541 a_7177_n1068.t3 a_7177_n1068.t4 298.839
R19542 a_7177_n1068.n0 a_7177_n1068.t5 280.405
R19543 a_7177_n1068.n1 a_7177_n1068.t0 200
R19544 a_7177_n1068.n1 a_7177_n1068.n0 172.311
R19545 a_7177_n1068.n2 a_7177_n1068.n1 24
R19546 a_7177_n1068.n1 a_7177_n1068.t1 21.212
R19547 a_4315_3184.t0 a_4315_3184.t1 242.857
R19548 a_372_211.n0 a_372_211.t2 358.166
R19549 a_372_211.t4 a_372_211.t3 337.399
R19550 a_372_211.t3 a_372_211.t5 285.986
R19551 a_372_211.n0 a_372_211.t4 282.573
R19552 a_372_211.n1 a_372_211.t1 202.857
R19553 a_372_211.n1 a_372_211.n0 173.817
R19554 a_372_211.n1 a_372_211.t0 20.826
R19555 a_372_211.n2 a_372_211.n1 20.689
R19556 a_277_196.n0 a_277_196.t2 362.857
R19557 a_277_196.t4 a_277_196.t3 337.399
R19558 a_277_196.t3 a_277_196.t5 298.839
R19559 a_277_196.n0 a_277_196.t4 280.405
R19560 a_277_196.n1 a_277_196.t0 200
R19561 a_277_196.n1 a_277_196.n0 172.311
R19562 a_277_196.n2 a_277_196.n1 24
R19563 a_277_196.n1 a_277_196.t1 21.212
R19564 a_553_n1770.n0 a_553_n1770.t1 160.619
R19565 a_553_n1770.t0 a_553_n1770.n0 151.153
R19566 SA_OUT[0].n1 SA_OUT[0].t3 661.027
R19567 SA_OUT[0].n1 SA_OUT[0].t4 392.255
R19568 SA_OUT[0].n2 SA_OUT[0].t2 223.716
R19569 SA_OUT[0].n0 SA_OUT[0].t0 153.977
R19570 SA_OUT[0].n2 SA_OUT[0].n1 143.764
R19571 SA_OUT[0].n0 SA_OUT[0].t1 59.86
R19572 SA_OUT[0] SA_OUT[0].n3 26.862
R19573 SA_OUT[0].n3 SA_OUT[0].n2 3.011
R19574 SA_OUT[0].n3 SA_OUT[0].n0 1.505
R19575 a_7067_3425.t0 a_7067_3425.t1 242.857
R19576 a_7039_n5850.n0 a_7039_n5850.t4 1465.51
R19577 a_7039_n5850.n0 a_7039_n5850.t3 712.44
R19578 a_7039_n5850.n1 a_7039_n5850.t0 375.067
R19579 a_7039_n5850.n1 a_7039_n5850.t1 272.668
R19580 a_7039_n5850.n2 a_7039_n5850.n0 143.764
R19581 a_7039_n5850.t2 a_7039_n5850.n2 78.193
R19582 a_7039_n5850.n2 a_7039_n5850.n1 4.517
R19583 ADC9_OUT[1].n0 ADC9_OUT[1].t4 1355.37
R19584 ADC9_OUT[1].n0 ADC9_OUT[1].t3 820.859
R19585 ADC9_OUT[1].n3 ADC9_OUT[1].t0 332.902
R19586 ADC9_OUT[1].n2 ADC9_OUT[1].t1 266.644
R19587 ADC9_OUT[1].n1 ADC9_OUT[1].n0 149.035
R19588 ADC9_OUT[1].n3 ADC9_OUT[1].n2 51.2
R19589 ADC9_OUT[1].n1 ADC9_OUT[1].t2 45.968
R19590 ADC9_OUT[1] ADC9_OUT[1].n3 45.927
R19591 ADC9_OUT[1].n2 ADC9_OUT[1].n1 17.317
R19592 a_5547_3907.n0 a_5547_3907.t1 358.166
R19593 a_5547_3907.t4 a_5547_3907.t5 337.399
R19594 a_5547_3907.t5 a_5547_3907.t3 285.986
R19595 a_5547_3907.n0 a_5547_3907.t4 282.573
R19596 a_5547_3907.n1 a_5547_3907.t0 202.857
R19597 a_5547_3907.n1 a_5547_3907.n0 173.817
R19598 a_5547_3907.n1 a_5547_3907.t2 20.826
R19599 a_5547_3907.n2 a_5547_3907.n1 20.689
R19600 a_3247_975.n0 a_3247_975.t2 358.166
R19601 a_3247_975.t4 a_3247_975.t5 337.399
R19602 a_3247_975.t5 a_3247_975.t3 285.986
R19603 a_3247_975.n0 a_3247_975.t4 282.573
R19604 a_3247_975.n1 a_3247_975.t0 202.857
R19605 a_3247_975.n1 a_3247_975.n0 173.817
R19606 a_3247_975.n1 a_3247_975.t1 20.826
R19607 a_3247_975.n2 a_3247_975.n1 20.689
R19608 a_352_n2234.n2 a_352_n2234.t0 282.97
R19609 a_352_n2234.n1 a_352_n2234.t2 240.683
R19610 a_352_n2234.n0 a_352_n2234.t3 209.208
R19611 a_352_n2234.n0 a_352_n2234.t4 194.167
R19612 a_352_n2234.t1 a_352_n2234.n2 183.404
R19613 a_352_n2234.n1 a_352_n2234.n0 14.805
R19614 a_352_n2234.n2 a_352_n2234.n1 6.415
R19615 a_277_n827.n0 a_277_n827.t1 362.857
R19616 a_277_n827.t3 a_277_n827.t4 337.399
R19617 a_277_n827.t4 a_277_n827.t5 298.839
R19618 a_277_n827.n0 a_277_n827.t3 280.405
R19619 a_277_n827.n1 a_277_n827.t0 200
R19620 a_277_n827.n1 a_277_n827.n0 172.311
R19621 a_277_n827.n2 a_277_n827.n1 24
R19622 a_277_n827.n1 a_277_n827.t2 21.212
R19623 a_372_n812.n0 a_372_n812.t2 358.166
R19624 a_372_n812.t3 a_372_n812.t5 337.399
R19625 a_372_n812.t5 a_372_n812.t4 285.986
R19626 a_372_n812.n0 a_372_n812.t3 282.573
R19627 a_372_n812.n1 a_372_n812.t0 202.857
R19628 a_372_n812.n1 a_372_n812.n0 173.817
R19629 a_372_n812.n1 a_372_n812.t1 20.826
R19630 a_372_n812.n2 a_372_n812.n1 20.689
R19631 a_7190_4445.t0 a_7190_4445.t1 242.857
R19632 a_1317_2421.t0 a_1317_2421.t1 242.857
R19633 a_6697_1698.n0 a_6697_1698.t2 358.166
R19634 a_6697_1698.t3 a_6697_1698.t4 337.399
R19635 a_6697_1698.t4 a_6697_1698.t5 285.986
R19636 a_6697_1698.n0 a_6697_1698.t3 282.573
R19637 a_6697_1698.n1 a_6697_1698.t0 202.857
R19638 a_6697_1698.n1 a_6697_1698.n0 173.817
R19639 a_6697_1698.n1 a_6697_1698.t1 20.826
R19640 a_6697_1698.n2 a_6697_1698.n1 20.689
R19641 a_1317_n271.t0 a_1317_n271.t1 242.857
R19642 a_742_n1053.t0 a_742_n1053.t1 242.857
R19643 a_1892_n812.t0 a_1892_n812.t1 242.857
R19644 a_3727_4671.n0 a_3727_4671.t2 362.857
R19645 a_3727_4671.t5 a_3727_4671.t3 337.399
R19646 a_3727_4671.t3 a_3727_4671.t4 298.839
R19647 a_3727_4671.n0 a_3727_4671.t5 280.405
R19648 a_3727_4671.n1 a_3727_4671.t0 200
R19649 a_3727_4671.n1 a_3727_4671.n0 172.311
R19650 a_3727_4671.n2 a_3727_4671.n1 24
R19651 a_3727_4671.n1 a_3727_4671.t1 21.212
R19652 a_8340_2180.t0 a_8340_2180.t1 242.857
R19653 a_947_3184.n0 a_947_3184.t1 358.166
R19654 a_947_3184.t5 a_947_3184.t3 337.399
R19655 a_947_3184.t3 a_947_3184.t4 285.986
R19656 a_947_3184.n0 a_947_3184.t5 282.573
R19657 a_947_3184.n1 a_947_3184.t0 202.857
R19658 a_947_3184.n1 a_947_3184.n0 173.817
R19659 a_947_3184.n1 a_947_3184.t2 20.826
R19660 a_947_3184.n2 a_947_3184.n1 20.689
R19661 a_852_3169.n0 a_852_3169.t1 362.857
R19662 a_852_3169.t3 a_852_3169.t4 337.399
R19663 a_852_3169.t4 a_852_3169.t5 298.839
R19664 a_852_3169.n0 a_852_3169.t3 280.405
R19665 a_852_3169.n1 a_852_3169.t2 200
R19666 a_852_3169.n1 a_852_3169.n0 172.311
R19667 a_852_3169.n2 a_852_3169.n1 24
R19668 a_852_3169.n1 a_852_3169.t0 21.212
R19669 a_3152_196.n0 a_3152_196.t0 362.857
R19670 a_3152_196.t4 a_3152_196.t3 337.399
R19671 a_3152_196.t3 a_3152_196.t5 298.839
R19672 a_3152_196.n0 a_3152_196.t4 280.405
R19673 a_3152_196.n1 a_3152_196.t1 200
R19674 a_3152_196.n1 a_3152_196.n0 172.311
R19675 a_3152_196.n2 a_3152_196.n1 24
R19676 a_3152_196.n1 a_3152_196.t2 21.212
R19677 a_3247_211.n0 a_3247_211.t1 358.166
R19678 a_3247_211.t5 a_3247_211.t4 337.399
R19679 a_3247_211.t4 a_3247_211.t3 285.986
R19680 a_3247_211.n0 a_3247_211.t5 282.573
R19681 a_3247_211.n1 a_3247_211.t2 202.857
R19682 a_3247_211.n1 a_3247_211.n0 173.817
R19683 a_3247_211.n1 a_3247_211.t0 20.826
R19684 a_3247_211.n2 a_3247_211.n1 20.689
R19685 a_1695_4887.n25 a_1695_4887.t27 561.971
R19686 a_1695_4887.n0 a_1695_4887.t5 449.944
R19687 a_1695_4887.t15 a_1695_4887.n25 108.636
R19688 a_1695_4887.n0 a_1695_4887.t6 74.821
R19689 a_1695_4887.n24 a_1695_4887.t22 63.519
R19690 a_1695_4887.n23 a_1695_4887.t1 63.519
R19691 a_1695_4887.n22 a_1695_4887.t14 63.519
R19692 a_1695_4887.n21 a_1695_4887.t16 63.519
R19693 a_1695_4887.n20 a_1695_4887.t13 63.519
R19694 a_1695_4887.n19 a_1695_4887.t19 63.519
R19695 a_1695_4887.n18 a_1695_4887.t20 63.519
R19696 a_1695_4887.n17 a_1695_4887.t10 63.519
R19697 a_1695_4887.n16 a_1695_4887.t4 63.519
R19698 a_1695_4887.n15 a_1695_4887.t8 63.519
R19699 a_1695_4887.n14 a_1695_4887.t23 63.519
R19700 a_1695_4887.n13 a_1695_4887.t21 63.519
R19701 a_1695_4887.n12 a_1695_4887.t18 63.519
R19702 a_1695_4887.n11 a_1695_4887.t11 63.519
R19703 a_1695_4887.n10 a_1695_4887.t12 63.519
R19704 a_1695_4887.n9 a_1695_4887.t24 63.519
R19705 a_1695_4887.n8 a_1695_4887.t0 63.519
R19706 a_1695_4887.n7 a_1695_4887.t3 63.519
R19707 a_1695_4887.n6 a_1695_4887.t2 63.519
R19708 a_1695_4887.n5 a_1695_4887.t26 63.519
R19709 a_1695_4887.n4 a_1695_4887.t9 63.519
R19710 a_1695_4887.n3 a_1695_4887.t17 63.519
R19711 a_1695_4887.n2 a_1695_4887.t25 63.519
R19712 a_1695_4887.n1 a_1695_4887.t7 63.519
R19713 a_1695_4887.n1 a_1695_4887.n0 8.619
R19714 a_1695_4887.n25 a_1695_4887.n24 2.946
R19715 a_1695_4887.n23 a_1695_4887.n22 2.524
R19716 a_1695_4887.n3 a_1695_4887.n2 2.498
R19717 a_1695_4887.n17 a_1695_4887.n16 2.364
R19718 a_1695_4887.n9 a_1695_4887.n8 2.355
R19719 a_1695_4887.n24 a_1695_4887.n23 1.998
R19720 a_1695_4887.n22 a_1695_4887.n21 1.998
R19721 a_1695_4887.n21 a_1695_4887.n20 1.998
R19722 a_1695_4887.n20 a_1695_4887.n19 1.998
R19723 a_1695_4887.n19 a_1695_4887.n18 1.998
R19724 a_1695_4887.n18 a_1695_4887.n17 1.998
R19725 a_1695_4887.n16 a_1695_4887.n15 1.998
R19726 a_1695_4887.n15 a_1695_4887.n14 1.998
R19727 a_1695_4887.n14 a_1695_4887.n13 1.998
R19728 a_1695_4887.n13 a_1695_4887.n12 1.998
R19729 a_1695_4887.n12 a_1695_4887.n11 1.998
R19730 a_1695_4887.n11 a_1695_4887.n10 1.998
R19731 a_1695_4887.n10 a_1695_4887.n9 1.998
R19732 a_1695_4887.n8 a_1695_4887.n7 1.998
R19733 a_1695_4887.n7 a_1695_4887.n6 1.998
R19734 a_1695_4887.n6 a_1695_4887.n5 1.998
R19735 a_1695_4887.n5 a_1695_4887.n4 1.998
R19736 a_1695_4887.n4 a_1695_4887.n3 1.998
R19737 a_1695_4887.n2 a_1695_4887.n1 1.998
R19738 a_1427_196.n0 a_1427_196.t1 362.857
R19739 a_1427_196.t4 a_1427_196.t3 337.399
R19740 a_1427_196.t3 a_1427_196.t5 298.839
R19741 a_1427_196.n0 a_1427_196.t4 280.405
R19742 a_1427_196.n1 a_1427_196.t2 200
R19743 a_1427_196.n1 a_1427_196.n0 172.311
R19744 a_1427_196.n2 a_1427_196.n1 24
R19745 a_1427_196.n1 a_1427_196.t0 21.212
R19746 a_2577_3892.n0 a_2577_3892.t2 362.857
R19747 a_2577_3892.t3 a_2577_3892.t4 337.399
R19748 a_2577_3892.t4 a_2577_3892.t5 298.839
R19749 a_2577_3892.n0 a_2577_3892.t3 280.405
R19750 a_2577_3892.n1 a_2577_3892.t0 200
R19751 a_2577_3892.n1 a_2577_3892.n0 172.311
R19752 a_2577_3892.n2 a_2577_3892.n1 24
R19753 a_2577_3892.n1 a_2577_3892.t1 21.212
R19754 a_2672_3907.n0 a_2672_3907.t2 358.166
R19755 a_2672_3907.t5 a_2672_3907.t3 337.399
R19756 a_2672_3907.t3 a_2672_3907.t4 285.986
R19757 a_2672_3907.n0 a_2672_3907.t5 282.573
R19758 a_2672_3907.n1 a_2672_3907.t0 202.857
R19759 a_2672_3907.n1 a_2672_3907.n0 173.817
R19760 a_2672_3907.n1 a_2672_3907.t1 20.826
R19761 a_2672_3907.n2 a_2672_3907.n1 20.689
R19762 a_852_2165.n0 a_852_2165.t2 362.857
R19763 a_852_2165.t4 a_852_2165.t5 337.399
R19764 a_852_2165.t5 a_852_2165.t3 298.839
R19765 a_852_2165.n0 a_852_2165.t4 280.405
R19766 a_852_2165.n1 a_852_2165.t0 200
R19767 a_852_2165.n1 a_852_2165.n0 172.311
R19768 a_852_2165.n2 a_852_2165.n1 24
R19769 a_852_2165.n1 a_852_2165.t1 21.212
R19770 a_865_2180.t0 a_865_2180.t1 242.857
R19771 a_6697_n812.n0 a_6697_n812.t1 358.166
R19772 a_6697_n812.t3 a_6697_n812.t4 337.399
R19773 a_6697_n812.t4 a_6697_n812.t5 285.986
R19774 a_6697_n812.n0 a_6697_n812.t3 282.573
R19775 a_6697_n812.n1 a_6697_n812.t0 202.857
R19776 a_6697_n812.n1 a_6697_n812.n0 173.817
R19777 a_6697_n812.n1 a_6697_n812.t2 20.826
R19778 a_6697_n812.n2 a_6697_n812.n1 20.689
R19779 a_6602_n827.n0 a_6602_n827.t2 362.857
R19780 a_6602_n827.t3 a_6602_n827.t5 337.399
R19781 a_6602_n827.t5 a_6602_n827.t4 298.839
R19782 a_6602_n827.n0 a_6602_n827.t3 280.405
R19783 a_6602_n827.n1 a_6602_n827.t0 200
R19784 a_6602_n827.n1 a_6602_n827.n0 172.311
R19785 a_6602_n827.n2 a_6602_n827.n1 24
R19786 a_6602_n827.n1 a_6602_n827.t1 21.212
R19787 a_3740_2943.t0 a_3740_2943.t1 242.857
R19788 a_3822_4445.n0 a_3822_4445.t0 358.166
R19789 a_3822_4445.t4 a_3822_4445.t3 337.399
R19790 a_3822_4445.t3 a_3822_4445.t5 285.986
R19791 a_3822_4445.n0 a_3822_4445.t4 282.573
R19792 a_3822_4445.n1 a_3822_4445.t2 202.857
R19793 a_3822_4445.n1 a_3822_4445.n0 173.817
R19794 a_3822_4445.n1 a_3822_4445.t1 20.826
R19795 a_3822_4445.n2 a_3822_4445.n1 20.689
R19796 a_3727_4430.n0 a_3727_4430.t1 362.857
R19797 a_3727_4430.t3 a_3727_4430.t4 337.399
R19798 a_3727_4430.t4 a_3727_4430.t5 298.839
R19799 a_3727_4430.n0 a_3727_4430.t3 280.405
R19800 a_3727_4430.n1 a_3727_4430.t2 200
R19801 a_3727_4430.n1 a_3727_4430.n0 172.311
R19802 a_3727_4430.n2 a_3727_4430.n1 24
R19803 a_3727_4430.n1 a_3727_4430.t0 21.212
R19804 a_4767_2180.t0 a_4767_2180.t1 242.857
R19805 a_2002_678.n0 a_2002_678.t0 362.857
R19806 a_2002_678.t5 a_2002_678.t4 337.399
R19807 a_2002_678.t4 a_2002_678.t3 298.839
R19808 a_2002_678.n0 a_2002_678.t5 280.405
R19809 a_2002_678.n1 a_2002_678.t2 200
R19810 a_2002_678.n1 a_2002_678.n0 172.311
R19811 a_2002_678.n2 a_2002_678.n1 24
R19812 a_2002_678.n1 a_2002_678.t1 21.212
R19813 a_2015_693.t0 a_2015_693.t1 242.857
R19814 a_3617_4148.t0 a_3617_4148.t1 242.857
R19815 a_277_1442.n0 a_277_1442.t2 362.857
R19816 a_277_1442.t3 a_277_1442.t4 337.399
R19817 a_277_1442.t4 a_277_1442.t5 298.839
R19818 a_277_1442.n0 a_277_1442.t3 280.405
R19819 a_277_1442.n1 a_277_1442.t0 200
R19820 a_277_1442.n1 a_277_1442.n0 172.311
R19821 a_277_1442.n2 a_277_1442.n1 24
R19822 a_277_1442.n1 a_277_1442.t1 21.212
R19823 a_867_n5092.t0 a_867_n5092.t1 42.705
R19824 a_902_n5293.n0 a_902_n5293.t0 65.063
R19825 a_902_n5293.n0 a_902_n5293.t2 42.011
R19826 a_902_n5293.t1 a_902_n5293.n0 2.113
R19827 Din[6].n0 Din[6].t1 215.292
R19828 Din[6].n0 Din[6].t0 187.376
R19829 Din[6] Din[6].n0 84.92
R19830 a_7272_1457.n0 a_7272_1457.t0 358.166
R19831 a_7272_1457.t3 a_7272_1457.t5 337.399
R19832 a_7272_1457.t5 a_7272_1457.t4 285.986
R19833 a_7272_1457.n0 a_7272_1457.t3 282.573
R19834 a_7272_1457.n1 a_7272_1457.t2 202.857
R19835 a_7272_1457.n1 a_7272_1457.n0 173.817
R19836 a_7272_1457.n1 a_7272_1457.t1 20.826
R19837 a_7272_1457.n2 a_7272_1457.n1 20.689
R19838 a_7177_1442.n0 a_7177_1442.t1 362.857
R19839 a_7177_1442.t3 a_7177_1442.t4 337.399
R19840 a_7177_1442.t4 a_7177_1442.t5 298.839
R19841 a_7177_1442.n0 a_7177_1442.t3 280.405
R19842 a_7177_1442.n1 a_7177_1442.t2 200
R19843 a_7177_1442.n1 a_7177_1442.n0 172.311
R19844 a_7177_1442.n2 a_7177_1442.n1 24
R19845 a_7177_1442.n1 a_7177_1442.t0 21.212
R19846 a_4877_196.n0 a_4877_196.t2 362.857
R19847 a_4877_196.t4 a_4877_196.t3 337.399
R19848 a_4877_196.t3 a_4877_196.t5 298.839
R19849 a_4877_196.n0 a_4877_196.t4 280.405
R19850 a_4877_196.n1 a_4877_196.t0 200
R19851 a_4877_196.n1 a_4877_196.n0 172.311
R19852 a_4877_196.n2 a_4877_196.n1 24
R19853 a_4877_196.n1 a_4877_196.t1 21.212
R19854 a_4972_211.n0 a_4972_211.t2 358.166
R19855 a_4972_211.t5 a_4972_211.t4 337.399
R19856 a_4972_211.t4 a_4972_211.t3 285.986
R19857 a_4972_211.n0 a_4972_211.t5 282.573
R19858 a_4972_211.n1 a_4972_211.t0 202.857
R19859 a_4972_211.n1 a_4972_211.n0 173.817
R19860 a_4972_211.n1 a_4972_211.t1 20.826
R19861 a_4972_211.n2 a_4972_211.n1 20.689
R19862 a_4767_452.t0 a_4767_452.t1 242.857
R19863 a_6602_4430.n0 a_6602_4430.t0 362.857
R19864 a_6602_4430.t3 a_6602_4430.t5 337.399
R19865 a_6602_4430.t5 a_6602_4430.t4 298.839
R19866 a_6602_4430.n0 a_6602_4430.t3 280.405
R19867 a_6602_4430.n1 a_6602_4430.t2 200
R19868 a_6602_4430.n1 a_6602_4430.n0 172.311
R19869 a_6602_4430.n2 a_6602_4430.n1 24
R19870 a_6602_4430.n1 a_6602_4430.t1 21.212
R19871 a_2590_2662.t0 a_2590_2662.t1 242.857
R19872 a_742_211.t0 a_742_211.t1 242.857
R19873 a_5547_n271.n0 a_5547_n271.t0 358.166
R19874 a_5547_n271.t4 a_5547_n271.t5 337.399
R19875 a_5547_n271.t5 a_5547_n271.t3 285.986
R19876 a_5547_n271.n0 a_5547_n271.t4 282.573
R19877 a_5547_n271.n1 a_5547_n271.t2 202.857
R19878 a_5547_n271.n1 a_5547_n271.n0 173.817
R19879 a_5547_n271.n1 a_5547_n271.t1 20.826
R19880 a_5547_n271.n2 a_5547_n271.n1 20.689
R19881 a_8488_n5293.t1 a_8488_n5293.t0 336.814
R19882 a_8429_n5338.t0 a_8429_n5338.t1 68.74
R19883 a_852_1683.n0 a_852_1683.t1 362.857
R19884 a_852_1683.t3 a_852_1683.t4 337.399
R19885 a_852_1683.t4 a_852_1683.t5 298.839
R19886 a_852_1683.n0 a_852_1683.t3 280.405
R19887 a_852_1683.n1 a_852_1683.t0 200
R19888 a_852_1683.n1 a_852_1683.n0 172.311
R19889 a_852_1683.n2 a_852_1683.n1 24
R19890 a_852_1683.n1 a_852_1683.t2 21.212
R19891 a_947_1698.n0 a_947_1698.t1 358.166
R19892 a_947_1698.t4 a_947_1698.t5 337.399
R19893 a_947_1698.t5 a_947_1698.t3 285.986
R19894 a_947_1698.n0 a_947_1698.t4 282.573
R19895 a_947_1698.n1 a_947_1698.t2 202.857
R19896 a_947_1698.n1 a_947_1698.n0 173.817
R19897 a_947_1698.n1 a_947_1698.t0 20.826
R19898 a_947_1698.n2 a_947_1698.n1 20.689
R19899 a_3740_693.t0 a_3740_693.t1 242.857
R19900 a_372_1457.n0 a_372_1457.t2 358.166
R19901 a_372_1457.t5 a_372_1457.t4 337.399
R19902 a_372_1457.t4 a_372_1457.t3 285.986
R19903 a_372_1457.n0 a_372_1457.t5 282.573
R19904 a_372_1457.n1 a_372_1457.t0 202.857
R19905 a_372_1457.n1 a_372_1457.n0 173.817
R19906 a_372_1457.n1 a_372_1457.t1 20.826
R19907 a_372_1457.n2 a_372_1457.n1 20.689
R19908 a_742_1457.t0 a_742_1457.t1 242.857
R19909 a_2311_n8583.n0 a_2311_n8583.t3 1465.51
R19910 a_2311_n8583.n0 a_2311_n8583.t4 712.44
R19911 a_2311_n8583.n1 a_2311_n8583.t0 375.067
R19912 a_2311_n8583.n1 a_2311_n8583.t2 272.668
R19913 a_2311_n8583.n2 a_2311_n8583.n0 143.764
R19914 a_2311_n8583.t1 a_2311_n8583.n2 78.193
R19915 a_2311_n8583.n2 a_2311_n8583.n1 4.517
R19916 ADC5_OUT[3].n0 ADC5_OUT[3].t3 1355.37
R19917 ADC5_OUT[3].n0 ADC5_OUT[3].t4 820.859
R19918 ADC5_OUT[3].n3 ADC5_OUT[3].t2 327.632
R19919 ADC5_OUT[3].n2 ADC5_OUT[3].t1 266.644
R19920 ADC5_OUT[3].n1 ADC5_OUT[3].n0 149.035
R19921 ADC5_OUT[3].n3 ADC5_OUT[3].n2 56.47
R19922 ADC5_OUT[3].n1 ADC5_OUT[3].t0 45.968
R19923 ADC5_OUT[3] ADC5_OUT[3].n3 22.24
R19924 ADC5_OUT[3].n2 ADC5_OUT[3].n1 17.317
R19925 a_2672_4445.n0 a_2672_4445.t1 358.166
R19926 a_2672_4445.t3 a_2672_4445.t4 337.399
R19927 a_2672_4445.t4 a_2672_4445.t5 285.986
R19928 a_2672_4445.n0 a_2672_4445.t3 282.573
R19929 a_2672_4445.n1 a_2672_4445.t2 202.857
R19930 a_2672_4445.n1 a_2672_4445.n0 173.817
R19931 a_2672_4445.n1 a_2672_4445.t0 20.826
R19932 a_2672_4445.n2 a_2672_4445.n1 20.689
R19933 a_2577_4430.n0 a_2577_4430.t1 362.857
R19934 a_2577_4430.t3 a_2577_4430.t4 337.399
R19935 a_2577_4430.t4 a_2577_4430.t5 298.839
R19936 a_2577_4430.n0 a_2577_4430.t3 280.405
R19937 a_2577_4430.n1 a_2577_4430.t2 200
R19938 a_2577_4430.n1 a_2577_4430.n0 172.311
R19939 a_2577_4430.n2 a_2577_4430.n1 24
R19940 a_2577_4430.n1 a_2577_4430.t0 21.212
R19941 a_277_3169.n0 a_277_3169.t2 362.857
R19942 a_277_3169.t5 a_277_3169.t3 337.399
R19943 a_277_3169.t3 a_277_3169.t4 298.839
R19944 a_277_3169.n0 a_277_3169.t5 280.405
R19945 a_277_3169.n1 a_277_3169.t0 200
R19946 a_277_3169.n1 a_277_3169.n0 172.311
R19947 a_277_3169.n2 a_277_3169.n1 24
R19948 a_277_3169.n1 a_277_3169.t1 21.212
R19949 a_372_3184.n0 a_372_3184.t2 358.166
R19950 a_372_3184.t3 a_372_3184.t5 337.399
R19951 a_372_3184.t5 a_372_3184.t4 285.986
R19952 a_372_3184.n0 a_372_3184.t3 282.573
R19953 a_372_3184.n1 a_372_3184.t0 202.857
R19954 a_372_3184.n1 a_372_3184.n0 173.817
R19955 a_372_3184.n1 a_372_3184.t1 20.826
R19956 a_372_3184.n2 a_372_3184.n1 20.689
R19957 ADC4_OUT[3].n0 ADC4_OUT[3].t4 1355.37
R19958 ADC4_OUT[3].n0 ADC4_OUT[3].t3 820.859
R19959 ADC4_OUT[3].n3 ADC4_OUT[3].t0 327.632
R19960 ADC4_OUT[3].n2 ADC4_OUT[3].t1 266.644
R19961 ADC4_OUT[3].n1 ADC4_OUT[3].n0 149.035
R19962 ADC4_OUT[3].n3 ADC4_OUT[3].n2 56.47
R19963 ADC4_OUT[3].n1 ADC4_OUT[3].t2 45.968
R19964 ADC4_OUT[3] ADC4_OUT[3].n3 22.187
R19965 ADC4_OUT[3].n2 ADC4_OUT[3].n1 17.317
R19966 a_1129_n8583.n0 a_1129_n8583.t4 1465.51
R19967 a_1129_n8583.n0 a_1129_n8583.t3 712.44
R19968 a_1129_n8583.n1 a_1129_n8583.t0 375.067
R19969 a_1129_n8583.n1 a_1129_n8583.t1 272.668
R19970 a_1129_n8583.n2 a_1129_n8583.n0 143.764
R19971 a_1129_n8583.t2 a_1129_n8583.n2 78.193
R19972 a_1129_n8583.n2 a_1129_n8583.n1 4.517
R19973 a_4972_n512.n0 a_4972_n512.t2 358.166
R19974 a_4972_n512.t3 a_4972_n512.t5 337.399
R19975 a_4972_n512.t5 a_4972_n512.t4 285.986
R19976 a_4972_n512.n0 a_4972_n512.t3 282.573
R19977 a_4972_n512.n1 a_4972_n512.t0 202.857
R19978 a_4972_n512.n1 a_4972_n512.n0 173.817
R19979 a_4972_n512.n1 a_4972_n512.t1 20.826
R19980 a_4972_n512.n2 a_4972_n512.n1 20.689
R19981 a_5547_3425.n0 a_5547_3425.t1 358.166
R19982 a_5547_3425.t4 a_5547_3425.t5 337.399
R19983 a_5547_3425.t5 a_5547_3425.t3 285.986
R19984 a_5547_3425.n0 a_5547_3425.t4 282.573
R19985 a_5547_3425.n1 a_5547_3425.t0 202.857
R19986 a_5547_3425.n1 a_5547_3425.n0 173.817
R19987 a_5547_3425.n1 a_5547_3425.t2 20.826
R19988 a_5547_3425.n2 a_5547_3425.n1 20.689
R19989 a_n2677_n4378.n3 a_n2677_n4378.t3 470.699
R19990 a_n2677_n4378.t4 a_n2677_n4378.t6 228.696
R19991 a_n2677_n4378.n2 a_n2677_n4378.t1 185.704
R19992 a_n2677_n4378.n3 a_n2677_n4378.n2 166.206
R19993 a_n2677_n4378.n0 a_n2677_n4378.t4 126.761
R19994 a_n2677_n4378.n1 a_n2677_n4378.t5 126.284
R19995 a_n2677_n4378.n1 a_n2677_n4378.t0 126.284
R19996 a_n2677_n4378.t2 a_n2677_n4378.n3 122.5
R19997 a_n2677_n4378.t0 a_n2677_n4378.n0 115.122
R19998 a_n2677_n4378.n0 a_n2677_n4378.t7 111.229
R19999 a_n2677_n4378.n2 a_n2677_n4378.n1 8.764
R20000 a_n2677_n6849.t0 a_n2677_n6849.t1 42.707
R20001 Din[11].n0 Din[11].t1 215.292
R20002 Din[11].n0 Din[11].t0 187.376
R20003 Din[11] Din[11].n0 84.92
R20004 a_3165_2421.t0 a_3165_2421.t1 242.857
R20005 a_6027_2406.n0 a_6027_2406.t2 362.857
R20006 a_6027_2406.t5 a_6027_2406.t3 337.399
R20007 a_6027_2406.t3 a_6027_2406.t4 298.839
R20008 a_6027_2406.n0 a_6027_2406.t5 280.405
R20009 a_6027_2406.n1 a_6027_2406.t0 200
R20010 a_6027_2406.n1 a_6027_2406.n0 172.311
R20011 a_6027_2406.n2 a_6027_2406.n1 24
R20012 a_6027_2406.n1 a_6027_2406.t1 21.212
R20013 a_6122_2421.n0 a_6122_2421.t1 358.166
R20014 a_6122_2421.t4 a_6122_2421.t3 337.399
R20015 a_6122_2421.t3 a_6122_2421.t5 285.986
R20016 a_6122_2421.n0 a_6122_2421.t4 282.573
R20017 a_6122_2421.n1 a_6122_2421.t2 202.857
R20018 a_6122_2421.n1 a_6122_2421.n0 173.817
R20019 a_6122_2421.n1 a_6122_2421.t0 20.826
R20020 a_6122_2421.n2 a_6122_2421.n1 20.689
R20021 a_6697_1216.n0 a_6697_1216.t1 358.166
R20022 a_6697_1216.t3 a_6697_1216.t4 337.399
R20023 a_6697_1216.t4 a_6697_1216.t5 285.986
R20024 a_6697_1216.n0 a_6697_1216.t3 282.573
R20025 a_6697_1216.n1 a_6697_1216.t2 202.857
R20026 a_6697_1216.n1 a_6697_1216.n0 173.817
R20027 a_6697_1216.n1 a_6697_1216.t0 20.826
R20028 a_6697_1216.n2 a_6697_1216.n1 20.689
R20029 a_7039_n7216.n0 a_7039_n7216.t4 1464.36
R20030 a_7039_n7216.n0 a_7039_n7216.t3 713.588
R20031 a_7039_n7216.n1 a_7039_n7216.t0 374.998
R20032 a_7039_n7216.n1 a_7039_n7216.t1 273.351
R20033 a_7039_n7216.n2 a_7039_n7216.n0 143.764
R20034 a_7039_n7216.t2 a_7039_n7216.n2 78.209
R20035 a_7039_n7216.n2 a_7039_n7216.n1 4.517
R20036 a_2097_693.n0 a_2097_693.t1 358.166
R20037 a_2097_693.t3 a_2097_693.t5 337.399
R20038 a_2097_693.t5 a_2097_693.t4 285.986
R20039 a_2097_693.n0 a_2097_693.t3 282.573
R20040 a_2097_693.n1 a_2097_693.t2 202.857
R20041 a_2097_693.n1 a_2097_693.n0 173.817
R20042 a_2097_693.n1 a_2097_693.t0 20.826
R20043 a_2097_693.n2 a_2097_693.n1 20.689
R20044 a_6027_n286.n0 a_6027_n286.t0 362.857
R20045 a_6027_n286.t5 a_6027_n286.t3 337.399
R20046 a_6027_n286.t3 a_6027_n286.t4 298.839
R20047 a_6027_n286.n0 a_6027_n286.t5 280.405
R20048 a_6027_n286.n1 a_6027_n286.t2 200
R20049 a_6027_n286.n1 a_6027_n286.n0 172.311
R20050 a_6027_n286.n2 a_6027_n286.n1 24
R20051 a_6027_n286.n1 a_6027_n286.t1 21.212
R20052 a_6122_n271.n0 a_6122_n271.t1 358.166
R20053 a_6122_n271.t3 a_6122_n271.t5 337.399
R20054 a_6122_n271.t5 a_6122_n271.t4 285.986
R20055 a_6122_n271.n0 a_6122_n271.t3 282.573
R20056 a_6122_n271.n1 a_6122_n271.t2 202.857
R20057 a_6122_n271.n1 a_6122_n271.n0 173.817
R20058 a_6122_n271.n1 a_6122_n271.t0 20.826
R20059 a_6122_n271.n2 a_6122_n271.n1 20.689
R20060 a_7272_4445.n0 a_7272_4445.t2 358.166
R20061 a_7272_4445.t4 a_7272_4445.t3 337.399
R20062 a_7272_4445.t3 a_7272_4445.t5 285.986
R20063 a_7272_4445.n0 a_7272_4445.t4 282.573
R20064 a_7272_4445.n1 a_7272_4445.t0 202.857
R20065 a_7272_4445.n1 a_7272_4445.n0 173.817
R20066 a_7272_4445.n1 a_7272_4445.t1 20.826
R20067 a_7272_4445.n2 a_7272_4445.n1 20.689
R20068 a_7177_4430.n0 a_7177_4430.t2 362.857
R20069 a_7177_4430.t5 a_7177_4430.t3 337.399
R20070 a_7177_4430.t3 a_7177_4430.t4 298.839
R20071 a_7177_4430.n0 a_7177_4430.t5 280.405
R20072 a_7177_4430.n1 a_7177_4430.t0 200
R20073 a_7177_4430.n1 a_7177_4430.n0 172.311
R20074 a_7177_4430.n2 a_7177_4430.n1 24
R20075 a_7177_4430.n1 a_7177_4430.t1 21.212
R20076 a_277_437.n0 a_277_437.t1 362.857
R20077 a_277_437.t3 a_277_437.t5 337.399
R20078 a_277_437.t5 a_277_437.t4 298.839
R20079 a_277_437.n0 a_277_437.t3 280.405
R20080 a_277_437.n1 a_277_437.t2 200
R20081 a_277_437.n1 a_277_437.n0 172.311
R20082 a_277_437.n2 a_277_437.n1 24
R20083 a_277_437.n1 a_277_437.t0 21.212
R20084 a_8068_n2086.t0 a_8068_n2086.t1 34.8
R20085 a_277_4133.n0 a_277_4133.t2 362.857
R20086 a_277_4133.t4 a_277_4133.t5 337.399
R20087 a_277_4133.t5 a_277_4133.t3 298.839
R20088 a_277_4133.n0 a_277_4133.t4 280.405
R20089 a_277_4133.n1 a_277_4133.t0 200
R20090 a_277_4133.n1 a_277_4133.n0 172.311
R20091 a_277_4133.n2 a_277_4133.n1 24
R20092 a_277_4133.n1 a_277_4133.t1 21.212
R20093 a_290_4148.t0 a_290_4148.t1 242.857
R20094 a_2672_3425.n0 a_2672_3425.t2 358.166
R20095 a_2672_3425.t5 a_2672_3425.t3 337.399
R20096 a_2672_3425.t3 a_2672_3425.t4 285.986
R20097 a_2672_3425.n0 a_2672_3425.t5 282.573
R20098 a_2672_3425.n1 a_2672_3425.t0 202.857
R20099 a_2672_3425.n1 a_2672_3425.n0 173.817
R20100 a_2672_3425.n1 a_2672_3425.t1 20.826
R20101 a_2672_3425.n2 a_2672_3425.n1 20.689
R20102 a_4192_4148.t0 a_4192_4148.t1 242.857
R20103 a_2381_n8071.n0 a_2381_n8071.t1 63.08
R20104 a_2381_n8071.t0 a_2381_n8071.n0 41.303
R20105 a_2381_n8071.n0 a_2381_n8071.t2 2.251
R20106 a_3247_693.n0 a_3247_693.t1 358.166
R20107 a_3247_693.t5 a_3247_693.t4 337.399
R20108 a_3247_693.t4 a_3247_693.t3 285.986
R20109 a_3247_693.n0 a_3247_693.t5 282.573
R20110 a_3247_693.n1 a_3247_693.t2 202.857
R20111 a_3247_693.n1 a_3247_693.n0 173.817
R20112 a_3247_693.n1 a_3247_693.t0 20.826
R20113 a_3247_693.n2 a_3247_693.n1 20.689
R20114 a_3617_693.t0 a_3617_693.t1 242.857
R20115 a_n2345_n8071.n0 a_n2345_n8071.t0 63.08
R20116 a_n2345_n8071.n0 a_n2345_n8071.t2 41.307
R20117 a_n2345_n8071.t1 a_n2345_n8071.n0 2.251
R20118 a_n2207_n8071.t0 a_n2207_n8071.t1 68.74
R20119 ADC7_OUT[3].n0 ADC7_OUT[3].t4 1355.37
R20120 ADC7_OUT[3].n0 ADC7_OUT[3].t3 820.859
R20121 ADC7_OUT[3].n3 ADC7_OUT[3].t0 332.902
R20122 ADC7_OUT[3].n2 ADC7_OUT[3].t2 266.644
R20123 ADC7_OUT[3].n1 ADC7_OUT[3].n0 149.035
R20124 ADC7_OUT[3].n3 ADC7_OUT[3].n2 51.2
R20125 ADC7_OUT[3].n1 ADC7_OUT[3].t1 45.968
R20126 ADC7_OUT[3] ADC7_OUT[3].n3 22.366
R20127 ADC7_OUT[3].n2 ADC7_OUT[3].n1 17.317
R20128 a_4302_3169.n0 a_4302_3169.t1 362.857
R20129 a_4302_3169.t3 a_4302_3169.t5 337.399
R20130 a_4302_3169.t5 a_4302_3169.t4 298.839
R20131 a_4302_3169.n0 a_4302_3169.t3 280.405
R20132 a_4302_3169.n1 a_4302_3169.t0 200
R20133 a_4302_3169.n1 a_4302_3169.n0 172.311
R20134 a_4302_3169.n2 a_4302_3169.n1 24
R20135 a_4302_3169.n1 a_4302_3169.t2 21.212
R20136 a_3235_n1770.n0 a_3235_n1770.t1 325.682
R20137 a_3235_n1770.t0 a_3235_n1770.n0 322.293
R20138 a_3235_n1770.n0 a_3235_n1770.t2 73.623
R20139 a_3277_n1770.t0 a_3277_n1770.n0 182.779
R20140 a_3277_n1770.n0 a_3277_n1770.t1 111.474
R20141 a_372_975.n0 a_372_975.t1 358.166
R20142 a_372_975.t3 a_372_975.t5 337.399
R20143 a_372_975.t5 a_372_975.t4 285.986
R20144 a_372_975.n0 a_372_975.t3 282.573
R20145 a_372_975.n1 a_372_975.t0 202.857
R20146 a_372_975.n1 a_372_975.n0 173.817
R20147 a_372_975.n1 a_372_975.t2 20.826
R20148 a_372_975.n2 a_372_975.n1 20.689
R20149 a_277_960.n0 a_277_960.t2 362.857
R20150 a_277_960.t3 a_277_960.t5 337.399
R20151 a_277_960.t5 a_277_960.t4 298.839
R20152 a_277_960.n0 a_277_960.t3 280.405
R20153 a_277_960.n1 a_277_960.t0 200
R20154 a_277_960.n1 a_277_960.n0 172.311
R20155 a_277_960.n2 a_277_960.n1 24
R20156 a_277_960.n1 a_277_960.t1 21.212
R20157 Din[8].n0 Din[8].t1 215.292
R20158 Din[8].n0 Din[8].t0 187.376
R20159 Din[8] Din[8].n0 84.911
R20160 a_5465_4148.t0 a_5465_4148.t1 242.857
R20161 a_8327_4133.n0 a_8327_4133.t2 362.857
R20162 a_8327_4133.t5 a_8327_4133.t3 337.399
R20163 a_8327_4133.t3 a_8327_4133.t4 298.839
R20164 a_8327_4133.n0 a_8327_4133.t5 280.405
R20165 a_8327_4133.n1 a_8327_4133.t0 200
R20166 a_8327_4133.n1 a_8327_4133.n0 172.311
R20167 a_8327_4133.n2 a_8327_4133.n1 24
R20168 a_8327_4133.n1 a_8327_4133.t1 21.212
R20169 a_8422_4148.n0 a_8422_4148.t2 358.166
R20170 a_8422_4148.t4 a_8422_4148.t3 337.399
R20171 a_8422_4148.t3 a_8422_4148.t5 285.986
R20172 a_8422_4148.n0 a_8422_4148.t4 282.573
R20173 a_8422_4148.n1 a_8422_4148.t0 202.857
R20174 a_8422_4148.n1 a_8422_4148.n0 173.817
R20175 a_8422_4148.n1 a_8422_4148.t1 20.826
R20176 a_8422_4148.n2 a_8422_4148.n1 20.689
R20177 a_8340_3184.t0 a_8340_3184.t1 242.857
R20178 a_5342_211.t0 a_5342_211.t1 242.857
R20179 a_13864_n8583.n0 a_13864_n8583.t4 1465.51
R20180 a_13864_n8583.n0 a_13864_n8583.t3 712.44
R20181 a_13864_n8583.n1 a_13864_n8583.t0 375.067
R20182 a_13864_n8583.n1 a_13864_n8583.t2 272.668
R20183 a_13864_n8583.n2 a_13864_n8583.n0 143.764
R20184 a_13864_n8583.t1 a_13864_n8583.n2 78.193
R20185 a_13864_n8583.n2 a_13864_n8583.n1 4.517
R20186 ADC15_OUT[3].n0 ADC15_OUT[3].t3 1355.37
R20187 ADC15_OUT[3].n0 ADC15_OUT[3].t4 820.859
R20188 ADC15_OUT[3].n3 ADC15_OUT[3].t0 336.667
R20189 ADC15_OUT[3].n2 ADC15_OUT[3].t1 266.644
R20190 ADC15_OUT[3].n1 ADC15_OUT[3].n0 149.035
R20191 ADC15_OUT[3].n3 ADC15_OUT[3].n2 47.435
R20192 ADC15_OUT[3].n1 ADC15_OUT[3].t2 45.968
R20193 ADC15_OUT[3] ADC15_OUT[3].n3 22.16
R20194 ADC15_OUT[3].n2 ADC15_OUT[3].n1 17.317
R20195 a_865_3184.t0 a_865_3184.t1 242.857
R20196 a_1427_2928.n0 a_1427_2928.t2 362.857
R20197 a_1427_2928.t5 a_1427_2928.t3 337.399
R20198 a_1427_2928.t3 a_1427_2928.t4 298.839
R20199 a_1427_2928.n0 a_1427_2928.t5 280.405
R20200 a_1427_2928.n1 a_1427_2928.t0 200
R20201 a_1427_2928.n1 a_1427_2928.n0 172.311
R20202 a_1427_2928.n2 a_1427_2928.n1 24
R20203 a_1427_2928.n1 a_1427_2928.t1 21.212
R20204 a_852_1201.n0 a_852_1201.t2 362.857
R20205 a_852_1201.t3 a_852_1201.t4 337.399
R20206 a_852_1201.t4 a_852_1201.t5 298.839
R20207 a_852_1201.n0 a_852_1201.t3 280.405
R20208 a_852_1201.n1 a_852_1201.t0 200
R20209 a_852_1201.n1 a_852_1201.n0 172.311
R20210 a_852_1201.n2 a_852_1201.n1 24
R20211 a_852_1201.n1 a_852_1201.t1 21.212
R20212 a_947_1216.n0 a_947_1216.t2 358.166
R20213 a_947_1216.t4 a_947_1216.t5 337.399
R20214 a_947_1216.t5 a_947_1216.t3 285.986
R20215 a_947_1216.n0 a_947_1216.t4 282.573
R20216 a_947_1216.n1 a_947_1216.t0 202.857
R20217 a_947_1216.n1 a_947_1216.n0 173.817
R20218 a_947_1216.n1 a_947_1216.t1 20.826
R20219 a_947_1216.n2 a_947_1216.n1 20.689
R20220 a_1129_n4483.n0 a_1129_n4483.t4 1464.36
R20221 a_1129_n4483.n0 a_1129_n4483.t3 713.588
R20222 a_1129_n4483.n1 a_1129_n4483.t0 374.998
R20223 a_1129_n4483.n1 a_1129_n4483.t2 273.351
R20224 a_1129_n4483.n2 a_1129_n4483.n0 143.764
R20225 a_1129_n4483.t1 a_1129_n4483.n2 78.209
R20226 a_1129_n4483.n2 a_1129_n4483.n1 4.517
R20227 a_2002_n1068.n0 a_2002_n1068.t0 362.857
R20228 a_2002_n1068.t4 a_2002_n1068.t5 337.399
R20229 a_2002_n1068.t5 a_2002_n1068.t3 298.839
R20230 a_2002_n1068.n0 a_2002_n1068.t4 280.405
R20231 a_2002_n1068.n1 a_2002_n1068.t2 200
R20232 a_2002_n1068.n1 a_2002_n1068.n0 172.311
R20233 a_2002_n1068.n2 a_2002_n1068.n1 24
R20234 a_2002_n1068.n1 a_2002_n1068.t1 21.212
R20235 a_2015_n1053.t0 a_2015_n1053.t1 242.857
R20236 a_7067_n812.t0 a_7067_n812.t1 242.857
R20237 a_5342_2421.t0 a_5342_2421.t1 242.857
R20238 a_7272_975.n0 a_7272_975.t1 358.166
R20239 a_7272_975.t3 a_7272_975.t5 337.399
R20240 a_7272_975.t5 a_7272_975.t4 285.986
R20241 a_7272_975.n0 a_7272_975.t3 282.573
R20242 a_7272_975.n1 a_7272_975.t0 202.857
R20243 a_7272_975.n1 a_7272_975.n0 173.817
R20244 a_7272_975.n1 a_7272_975.t2 20.826
R20245 a_7272_975.n2 a_7272_975.n1 20.689
R20246 a_852_n827.n0 a_852_n827.t1 362.857
R20247 a_852_n827.t3 a_852_n827.t4 337.399
R20248 a_852_n827.t4 a_852_n827.t5 298.839
R20249 a_852_n827.n0 a_852_n827.t3 280.405
R20250 a_852_n827.n1 a_852_n827.t0 200
R20251 a_852_n827.n1 a_852_n827.n0 172.311
R20252 a_852_n827.n2 a_852_n827.n1 24
R20253 a_852_n827.n1 a_852_n827.t2 21.212
R20254 a_4397_3184.n0 a_4397_3184.t2 358.166
R20255 a_4397_3184.t4 a_4397_3184.t5 337.399
R20256 a_4397_3184.t5 a_4397_3184.t3 285.986
R20257 a_4397_3184.n0 a_4397_3184.t4 282.573
R20258 a_4397_3184.n1 a_4397_3184.t0 202.857
R20259 a_4397_3184.n1 a_4397_3184.n0 173.817
R20260 a_4397_3184.n1 a_4397_3184.t1 20.826
R20261 a_4397_3184.n2 a_4397_3184.n1 20.689
R20262 a_4767_3184.t0 a_4767_3184.t1 242.857
R20263 a_5342_n271.t0 a_5342_n271.t1 242.857
R20264 a_5452_3892.n0 a_5452_3892.t2 362.857
R20265 a_5452_3892.t4 a_5452_3892.t5 337.399
R20266 a_5452_3892.t5 a_5452_3892.t3 298.839
R20267 a_5452_3892.n0 a_5452_3892.t4 280.405
R20268 a_5452_3892.n1 a_5452_3892.t0 200
R20269 a_5452_3892.n1 a_5452_3892.n0 172.311
R20270 a_5452_3892.n2 a_5452_3892.n1 24
R20271 a_5452_3892.n1 a_5452_3892.t1 21.212
R20272 a_5465_3907.t0 a_5465_3907.t1 242.857
R20273 a_2672_2662.n0 a_2672_2662.t2 358.166
R20274 a_2672_2662.t5 a_2672_2662.t3 337.399
R20275 a_2672_2662.t3 a_2672_2662.t4 285.986
R20276 a_2672_2662.n0 a_2672_2662.t5 282.573
R20277 a_2672_2662.n1 a_2672_2662.t0 202.857
R20278 a_2672_2662.n1 a_2672_2662.n0 173.817
R20279 a_2672_2662.n1 a_2672_2662.t1 20.826
R20280 a_2672_2662.n2 a_2672_2662.n1 20.689
R20281 a_2577_2647.n0 a_2577_2647.t1 362.857
R20282 a_2577_2647.t5 a_2577_2647.t3 337.399
R20283 a_2577_2647.t3 a_2577_2647.t4 298.839
R20284 a_2577_2647.n0 a_2577_2647.t5 280.405
R20285 a_2577_2647.n1 a_2577_2647.t2 200
R20286 a_2577_2647.n1 a_2577_2647.n0 172.311
R20287 a_2577_2647.n2 a_2577_2647.n1 24
R20288 a_2577_2647.n1 a_2577_2647.t0 21.212
R20289 a_6615_2421.t0 a_6615_2421.t1 242.857
R20290 ADC2_OUT[3].n0 ADC2_OUT[3].t4 1355.37
R20291 ADC2_OUT[3].n0 ADC2_OUT[3].t3 820.859
R20292 ADC2_OUT[3].n3 ADC2_OUT[3].t0 326.126
R20293 ADC2_OUT[3].n2 ADC2_OUT[3].t1 266.644
R20294 ADC2_OUT[3].n1 ADC2_OUT[3].n0 149.035
R20295 ADC2_OUT[3].n3 ADC2_OUT[3].n2 57.976
R20296 ADC2_OUT[3].n1 ADC2_OUT[3].t2 45.968
R20297 ADC2_OUT[3] ADC2_OUT[3].n3 22.079
R20298 ADC2_OUT[3].n2 ADC2_OUT[3].n1 17.317
R20299 a_10362_n3770.n0 a_10362_n3770.t0 65.064
R20300 a_10362_n3770.n0 a_10362_n3770.t2 42.011
R20301 a_10362_n3770.t1 a_10362_n3770.n0 2.113
R20302 a_8985_n1770.n0 a_8985_n1770.t1 325.682
R20303 a_8985_n1770.n0 a_8985_n1770.t2 322.294
R20304 a_8985_n1770.t0 a_8985_n1770.n0 73.623
R20305 a_1533_n953.n25 a_1533_n953.t27 561.971
R20306 a_1533_n953.n0 a_1533_n953.t6 461.908
R20307 a_1533_n953.t15 a_1533_n953.n25 108.635
R20308 a_1533_n953.n0 a_1533_n953.t5 79.512
R20309 a_1533_n953.n24 a_1533_n953.t22 65.401
R20310 a_1533_n953.n23 a_1533_n953.t1 65.401
R20311 a_1533_n953.n22 a_1533_n953.t14 65.401
R20312 a_1533_n953.n21 a_1533_n953.t16 65.401
R20313 a_1533_n953.n20 a_1533_n953.t13 65.401
R20314 a_1533_n953.n19 a_1533_n953.t19 65.401
R20315 a_1533_n953.n18 a_1533_n953.t20 65.401
R20316 a_1533_n953.n17 a_1533_n953.t10 65.401
R20317 a_1533_n953.n16 a_1533_n953.t4 65.401
R20318 a_1533_n953.n15 a_1533_n953.t8 65.401
R20319 a_1533_n953.n14 a_1533_n953.t23 65.401
R20320 a_1533_n953.n13 a_1533_n953.t21 65.401
R20321 a_1533_n953.n12 a_1533_n953.t18 65.401
R20322 a_1533_n953.n11 a_1533_n953.t11 65.401
R20323 a_1533_n953.n10 a_1533_n953.t12 65.401
R20324 a_1533_n953.n9 a_1533_n953.t24 65.401
R20325 a_1533_n953.n8 a_1533_n953.t0 65.401
R20326 a_1533_n953.n7 a_1533_n953.t3 65.401
R20327 a_1533_n953.n6 a_1533_n953.t2 65.401
R20328 a_1533_n953.n5 a_1533_n953.t26 65.401
R20329 a_1533_n953.n4 a_1533_n953.t9 65.401
R20330 a_1533_n953.n3 a_1533_n953.t17 65.401
R20331 a_1533_n953.n2 a_1533_n953.t25 65.401
R20332 a_1533_n953.n1 a_1533_n953.t7 65.401
R20333 a_1533_n953.n1 a_1533_n953.n0 5.64
R20334 a_1533_n953.n25 a_1533_n953.n24 4.438
R20335 a_1533_n953.n23 a_1533_n953.n22 2.524
R20336 a_1533_n953.n3 a_1533_n953.n2 2.498
R20337 a_1533_n953.n17 a_1533_n953.n16 2.364
R20338 a_1533_n953.n9 a_1533_n953.n8 2.355
R20339 a_1533_n953.n2 a_1533_n953.n1 1.998
R20340 a_1533_n953.n4 a_1533_n953.n3 1.998
R20341 a_1533_n953.n5 a_1533_n953.n4 1.998
R20342 a_1533_n953.n6 a_1533_n953.n5 1.998
R20343 a_1533_n953.n7 a_1533_n953.n6 1.998
R20344 a_1533_n953.n8 a_1533_n953.n7 1.998
R20345 a_1533_n953.n10 a_1533_n953.n9 1.998
R20346 a_1533_n953.n11 a_1533_n953.n10 1.998
R20347 a_1533_n953.n12 a_1533_n953.n11 1.998
R20348 a_1533_n953.n13 a_1533_n953.n12 1.998
R20349 a_1533_n953.n14 a_1533_n953.n13 1.998
R20350 a_1533_n953.n15 a_1533_n953.n14 1.998
R20351 a_1533_n953.n16 a_1533_n953.n15 1.998
R20352 a_1533_n953.n18 a_1533_n953.n17 1.998
R20353 a_1533_n953.n19 a_1533_n953.n18 1.998
R20354 a_1533_n953.n20 a_1533_n953.n19 1.998
R20355 a_1533_n953.n21 a_1533_n953.n20 1.998
R20356 a_1533_n953.n22 a_1533_n953.n21 1.998
R20357 a_1533_n953.n24 a_1533_n953.n23 1.998
R20358 a_1510_n1770.n0 a_1510_n1770.t2 322.294
R20359 a_1510_n1770.n1 a_1510_n1770.n0 229.466
R20360 a_1510_n1770.t0 a_1510_n1770.n1 151.15
R20361 a_1510_n1770.n0 a_1510_n1770.t1 73.623
R20362 a_1552_n1770.t0 a_1552_n1770.n0 182.779
R20363 a_1552_n1770.n0 a_1552_n1770.t1 111.474
R20364 a_2577_1924.n0 a_2577_1924.t1 362.857
R20365 a_2577_1924.t4 a_2577_1924.t5 337.399
R20366 a_2577_1924.t5 a_2577_1924.t3 298.839
R20367 a_2577_1924.n0 a_2577_1924.t4 280.405
R20368 a_2577_1924.n1 a_2577_1924.t0 200
R20369 a_2577_1924.n1 a_2577_1924.n0 172.311
R20370 a_2577_1924.n2 a_2577_1924.n1 24
R20371 a_2577_1924.n1 a_2577_1924.t2 21.212
R20372 a_2590_1939.t0 a_2590_1939.t1 242.857
R20373 a_277_4671.n0 a_277_4671.t0 362.857
R20374 a_277_4671.t3 a_277_4671.t4 337.399
R20375 a_277_4671.t4 a_277_4671.t5 298.839
R20376 a_277_4671.n0 a_277_4671.t3 280.405
R20377 a_277_4671.n1 a_277_4671.t1 200
R20378 a_277_4671.n1 a_277_4671.n0 172.311
R20379 a_277_4671.n2 a_277_4671.n1 24
R20380 a_277_4671.n1 a_277_4671.t2 21.212
R20381 a_7752_2928.n0 a_7752_2928.t2 362.857
R20382 a_7752_2928.t4 a_7752_2928.t5 337.399
R20383 a_7752_2928.t5 a_7752_2928.t3 298.839
R20384 a_7752_2928.n0 a_7752_2928.t4 280.405
R20385 a_7752_2928.n1 a_7752_2928.t0 200
R20386 a_7752_2928.n1 a_7752_2928.n0 172.311
R20387 a_7752_2928.n2 a_7752_2928.n1 24
R20388 a_7752_2928.n1 a_7752_2928.t1 21.212
R20389 a_7765_2943.t0 a_7765_2943.t1 242.857
R20390 a_7272_4686.n0 a_7272_4686.t1 358.166
R20391 a_7272_4686.t3 a_7272_4686.t5 337.399
R20392 a_7272_4686.t5 a_7272_4686.t4 285.986
R20393 a_7272_4686.n0 a_7272_4686.t3 282.573
R20394 a_7272_4686.n1 a_7272_4686.t0 202.857
R20395 a_7272_4686.n1 a_7272_4686.n0 173.817
R20396 a_7272_4686.n1 a_7272_4686.t2 20.826
R20397 a_7272_4686.n2 a_7272_4686.n1 20.689
R20398 a_7177_4671.n0 a_7177_4671.t2 362.857
R20399 a_7177_4671.t3 a_7177_4671.t4 337.399
R20400 a_7177_4671.t4 a_7177_4671.t5 298.839
R20401 a_7177_4671.n0 a_7177_4671.t3 280.405
R20402 a_7177_4671.n1 a_7177_4671.t0 200
R20403 a_7177_4671.n1 a_7177_4671.n0 172.311
R20404 a_7177_4671.n2 a_7177_4671.n1 24
R20405 a_7177_4671.n1 a_7177_4671.t1 21.212
R20406 Din[13].n0 Din[13].t1 215.292
R20407 Din[13].n0 Din[13].t0 187.376
R20408 Din[13] Din[13].n0 84.912
R20409 a_7642_4148.t0 a_7642_4148.t1 242.857
R20410 a_8792_2180.t0 a_8792_2180.t1 242.857
R20411 a_2577_2165.n0 a_2577_2165.t2 362.857
R20412 a_2577_2165.t3 a_2577_2165.t4 337.399
R20413 a_2577_2165.t4 a_2577_2165.t5 298.839
R20414 a_2577_2165.n0 a_2577_2165.t3 280.405
R20415 a_2577_2165.n1 a_2577_2165.t0 200
R20416 a_2577_2165.n1 a_2577_2165.n0 172.311
R20417 a_2577_2165.n2 a_2577_2165.n1 24
R20418 a_2577_2165.n1 a_2577_2165.t1 21.212
R20419 a_372_1698.n0 a_372_1698.t2 358.166
R20420 a_372_1698.t3 a_372_1698.t5 337.399
R20421 a_372_1698.t5 a_372_1698.t4 285.986
R20422 a_372_1698.n0 a_372_1698.t3 282.573
R20423 a_372_1698.n1 a_372_1698.t1 202.857
R20424 a_372_1698.n1 a_372_1698.n0 173.817
R20425 a_372_1698.n1 a_372_1698.t0 20.826
R20426 a_372_1698.n2 a_372_1698.n1 20.689
R20427 a_n3792_n6503.n0 a_n3792_n6503.t0 65.064
R20428 a_n3792_n6503.n0 a_n3792_n6503.t2 42.011
R20429 a_n3792_n6503.t1 a_n3792_n6503.n0 2.113
R20430 a_9218_n2086.t0 a_9218_n2086.t1 34.8
R20431 a_1427_4133.n0 a_1427_4133.t1 362.857
R20432 a_1427_4133.t3 a_1427_4133.t4 337.399
R20433 a_1427_4133.t4 a_1427_4133.t5 298.839
R20434 a_1427_4133.n0 a_1427_4133.t3 280.405
R20435 a_1427_4133.n1 a_1427_4133.t0 200
R20436 a_1427_4133.n1 a_1427_4133.n0 172.311
R20437 a_1427_4133.n2 a_1427_4133.n1 24
R20438 a_1427_4133.n1 a_1427_4133.t2 21.212
R20439 a_8915_4148.t0 a_8915_4148.t1 242.857
R20440 a_3247_2421.n0 a_3247_2421.t2 358.166
R20441 a_3247_2421.t5 a_3247_2421.t3 337.399
R20442 a_3247_2421.t3 a_3247_2421.t4 285.986
R20443 a_3247_2421.n0 a_3247_2421.t5 282.573
R20444 a_3247_2421.n1 a_3247_2421.t0 202.857
R20445 a_3247_2421.n1 a_3247_2421.n0 173.817
R20446 a_3247_2421.n1 a_3247_2421.t1 20.826
R20447 a_3247_2421.n2 a_3247_2421.n1 20.689
R20448 a_3152_2406.n0 a_3152_2406.t1 362.857
R20449 a_3152_2406.t3 a_3152_2406.t4 337.399
R20450 a_3152_2406.t4 a_3152_2406.t5 298.839
R20451 a_3152_2406.n0 a_3152_2406.t3 280.405
R20452 a_3152_2406.n1 a_3152_2406.t2 200
R20453 a_3152_2406.n1 a_3152_2406.n0 172.311
R20454 a_3152_2406.n2 a_3152_2406.n1 24
R20455 a_3152_2406.n1 a_3152_2406.t0 21.212
R20456 ADC14_OUT[1].n0 ADC14_OUT[1].t4 1355.37
R20457 ADC14_OUT[1].n0 ADC14_OUT[1].t3 820.859
R20458 ADC14_OUT[1].n3 ADC14_OUT[1].t0 317.091
R20459 ADC14_OUT[1].n2 ADC14_OUT[1].t1 266.644
R20460 ADC14_OUT[1].n1 ADC14_OUT[1].n0 149.035
R20461 ADC14_OUT[1].n3 ADC14_OUT[1].n2 67.011
R20462 ADC14_OUT[1] ADC14_OUT[1].n3 45.99
R20463 ADC14_OUT[1].n1 ADC14_OUT[1].t2 45.968
R20464 ADC14_OUT[1].n2 ADC14_OUT[1].n1 17.317
R20465 a_12963_n5850.n0 a_12963_n5850.t4 1465.51
R20466 a_12963_n5850.n0 a_12963_n5850.t3 712.44
R20467 a_12963_n5850.n1 a_12963_n5850.t0 375.067
R20468 a_12963_n5850.n1 a_12963_n5850.t1 272.668
R20469 a_12963_n5850.n2 a_12963_n5850.n0 143.764
R20470 a_12963_n5850.t2 a_12963_n5850.n2 78.193
R20471 a_12963_n5850.n2 a_12963_n5850.n1 4.517
R20472 a_372_4686.n0 a_372_4686.t1 358.166
R20473 a_372_4686.t5 a_372_4686.t4 337.399
R20474 a_372_4686.t4 a_372_4686.t3 285.986
R20475 a_372_4686.n0 a_372_4686.t5 282.573
R20476 a_372_4686.n1 a_372_4686.t2 202.857
R20477 a_372_4686.n1 a_372_4686.n0 173.817
R20478 a_372_4686.n1 a_372_4686.t0 20.826
R20479 a_372_4686.n2 a_372_4686.n1 20.689
R20480 a_742_4686.t0 a_742_4686.t1 242.857
R20481 a_n314_n6849.t0 a_n314_n6849.t1 42.707
R20482 a_4890_3666.t0 a_4890_3666.t1 242.857
R20483 a_7272_n30.n0 a_7272_n30.t1 358.166
R20484 a_7272_n30.t4 a_7272_n30.t5 337.399
R20485 a_7272_n30.t5 a_7272_n30.t3 285.986
R20486 a_7272_n30.n0 a_7272_n30.t4 282.573
R20487 a_7272_n30.n1 a_7272_n30.t2 202.857
R20488 a_7272_n30.n1 a_7272_n30.n0 173.817
R20489 a_7272_n30.n1 a_7272_n30.t0 20.826
R20490 a_7272_n30.n2 a_7272_n30.n1 20.689
R20491 a_8291_n7203.n0 a_8291_n7203.t1 63.08
R20492 a_8291_n7203.t0 a_8291_n7203.n0 41.306
R20493 a_8291_n7203.n0 a_8291_n7203.t2 2.251
R20494 a_4385_n1770.n0 a_4385_n1770.t1 325.682
R20495 a_4385_n1770.n0 a_4385_n1770.t2 322.294
R20496 a_4385_n1770.t0 a_4385_n1770.n0 73.623
R20497 a_4427_n1770.t0 a_4427_n1770.t1 213.924
R20498 Din[14].n0 Din[14].t0 215.292
R20499 Din[14].n0 Din[14].t1 187.376
R20500 Din[14] Din[14].n0 84.947
R20501 a_8402_n2234.n2 a_8402_n2234.t1 282.97
R20502 a_8402_n2234.n1 a_8402_n2234.t4 240.683
R20503 a_8402_n2234.n0 a_8402_n2234.t2 209.208
R20504 a_8402_n2234.n0 a_8402_n2234.t3 194.167
R20505 a_8402_n2234.t0 a_8402_n2234.n2 183.404
R20506 a_8402_n2234.n1 a_8402_n2234.n0 14.805
R20507 a_8402_n2234.n2 a_8402_n2234.n1 6.415
R20508 a_6697_4445.n0 a_6697_4445.t1 358.166
R20509 a_6697_4445.t3 a_6697_4445.t4 337.399
R20510 a_6697_4445.t4 a_6697_4445.t5 285.986
R20511 a_6697_4445.n0 a_6697_4445.t3 282.573
R20512 a_6697_4445.n1 a_6697_4445.t2 202.857
R20513 a_6697_4445.n1 a_6697_4445.n0 173.817
R20514 a_6697_4445.n1 a_6697_4445.t0 20.826
R20515 a_6697_4445.n2 a_6697_4445.n1 20.689
R20516 a_6122_n30.n0 a_6122_n30.t2 358.166
R20517 a_6122_n30.t4 a_6122_n30.t5 337.399
R20518 a_6122_n30.t5 a_6122_n30.t3 285.986
R20519 a_6122_n30.n0 a_6122_n30.t4 282.573
R20520 a_6122_n30.n1 a_6122_n30.t0 202.857
R20521 a_6122_n30.n1 a_6122_n30.n0 173.817
R20522 a_6122_n30.n1 a_6122_n30.t1 20.826
R20523 a_6122_n30.n2 a_6122_n30.n1 20.689
R20524 a_6492_n30.t0 a_6492_n30.t1 242.857
R20525 a_8902_3892.n0 a_8902_3892.t1 362.857
R20526 a_8902_3892.t5 a_8902_3892.t4 337.399
R20527 a_8902_3892.t4 a_8902_3892.t3 298.839
R20528 a_8902_3892.n0 a_8902_3892.t5 280.405
R20529 a_8902_3892.n1 a_8902_3892.t0 200
R20530 a_8902_3892.n1 a_8902_3892.n0 172.311
R20531 a_8902_3892.n2 a_8902_3892.n1 24
R20532 a_8902_3892.n1 a_8902_3892.t2 21.212
R20533 a_8915_3907.t0 a_8915_3907.t1 242.857
R20534 a_5547_4148.n0 a_5547_4148.t0 358.166
R20535 a_5547_4148.t5 a_5547_4148.t3 337.399
R20536 a_5547_4148.t3 a_5547_4148.t4 285.986
R20537 a_5547_4148.n0 a_5547_4148.t5 282.573
R20538 a_5547_4148.n1 a_5547_4148.t2 202.857
R20539 a_5547_4148.n1 a_5547_4148.n0 173.817
R20540 a_5547_4148.n1 a_5547_4148.t1 20.826
R20541 a_5547_4148.n2 a_5547_4148.n1 20.689
R20542 a_5452_4133.n0 a_5452_4133.t1 362.857
R20543 a_5452_4133.t3 a_5452_4133.t4 337.399
R20544 a_5452_4133.t4 a_5452_4133.t5 298.839
R20545 a_5452_4133.n0 a_5452_4133.t3 280.405
R20546 a_5452_4133.n1 a_5452_4133.t2 200
R20547 a_5452_4133.n1 a_5452_4133.n0 172.311
R20548 a_5452_4133.n2 a_5452_4133.n1 24
R20549 a_5452_4133.n1 a_5452_4133.t0 21.212
R20550 a_5452_3410.n0 a_5452_3410.t2 362.857
R20551 a_5452_3410.t4 a_5452_3410.t5 337.399
R20552 a_5452_3410.t5 a_5452_3410.t3 298.839
R20553 a_5452_3410.n0 a_5452_3410.t4 280.405
R20554 a_5452_3410.n1 a_5452_3410.t0 200
R20555 a_5452_3410.n1 a_5452_3410.n0 172.311
R20556 a_5452_3410.n2 a_5452_3410.n1 24
R20557 a_5452_3410.n1 a_5452_3410.t1 21.212
R20558 a_5465_3425.t0 a_5465_3425.t1 242.857
R20559 a_7190_2421.t0 a_7190_2421.t1 242.857
R20560 a_3247_1939.n0 a_3247_1939.t1 358.166
R20561 a_3247_1939.t4 a_3247_1939.t5 337.399
R20562 a_3247_1939.t5 a_3247_1939.t3 285.986
R20563 a_3247_1939.n0 a_3247_1939.t4 282.573
R20564 a_3247_1939.n1 a_3247_1939.t2 202.857
R20565 a_3247_1939.n1 a_3247_1939.n0 173.817
R20566 a_3247_1939.n1 a_3247_1939.t0 20.826
R20567 a_3247_1939.n2 a_3247_1939.n1 20.689
R20568 a_3617_1939.t0 a_3617_1939.t1 242.857
R20569 a_3727_2647.n0 a_3727_2647.t1 362.857
R20570 a_3727_2647.t5 a_3727_2647.t3 337.399
R20571 a_3727_2647.t3 a_3727_2647.t4 298.839
R20572 a_3727_2647.n0 a_3727_2647.t5 280.405
R20573 a_3727_2647.n1 a_3727_2647.t2 200
R20574 a_3727_2647.n1 a_3727_2647.n0 172.311
R20575 a_3727_2647.n2 a_3727_2647.n1 24
R20576 a_3727_2647.n1 a_3727_2647.t0 21.212
R20577 a_7642_n30.t0 a_7642_n30.t1 242.857
R20578 a_9367_n512.t0 a_9367_n512.t1 242.857
R20579 a_3231_n5092.t0 a_3231_n5092.t1 42.705
R20580 a_3266_n5293.n0 a_3266_n5293.t0 65.064
R20581 a_3266_n5293.t1 a_3266_n5293.n0 42.011
R20582 a_3266_n5293.n0 a_3266_n5293.t2 2.113
R20583 a_3822_2421.n0 a_3822_2421.t0 358.166
R20584 a_3822_2421.t4 a_3822_2421.t3 337.399
R20585 a_3822_2421.t3 a_3822_2421.t5 285.986
R20586 a_3822_2421.n0 a_3822_2421.t4 282.573
R20587 a_3822_2421.n1 a_3822_2421.t2 202.857
R20588 a_3822_2421.n1 a_3822_2421.n0 173.817
R20589 a_3822_2421.n1 a_3822_2421.t1 20.826
R20590 a_3822_2421.n2 a_3822_2421.n1 20.689
R20591 a_3727_2406.n0 a_3727_2406.t1 362.857
R20592 a_3727_2406.t3 a_3727_2406.t4 337.399
R20593 a_3727_2406.t4 a_3727_2406.t5 298.839
R20594 a_3727_2406.n0 a_3727_2406.t3 280.405
R20595 a_3727_2406.n1 a_3727_2406.t2 200
R20596 a_3727_2406.n1 a_3727_2406.n0 172.311
R20597 a_3727_2406.n2 a_3727_2406.n1 24
R20598 a_3727_2406.n1 a_3727_2406.t0 21.212
R20599 a_3822_1457.n0 a_3822_1457.t1 358.166
R20600 a_3822_1457.t5 a_3822_1457.t4 337.399
R20601 a_3822_1457.t4 a_3822_1457.t3 285.986
R20602 a_3822_1457.n0 a_3822_1457.t5 282.573
R20603 a_3822_1457.n1 a_3822_1457.t2 202.857
R20604 a_3822_1457.n1 a_3822_1457.n0 173.817
R20605 a_3822_1457.n1 a_3822_1457.t0 20.826
R20606 a_3822_1457.n2 a_3822_1457.n1 20.689
R20607 a_5452_960.n0 a_5452_960.t1 362.857
R20608 a_5452_960.t4 a_5452_960.t3 337.399
R20609 a_5452_960.t3 a_5452_960.t5 298.839
R20610 a_5452_960.n0 a_5452_960.t4 280.405
R20611 a_5452_960.n1 a_5452_960.t0 200
R20612 a_5452_960.n1 a_5452_960.n0 172.311
R20613 a_5452_960.n2 a_5452_960.n1 24
R20614 a_5452_960.n1 a_5452_960.t2 21.212
R20615 a_5547_975.n0 a_5547_975.t2 358.166
R20616 a_5547_975.t4 a_5547_975.t5 337.399
R20617 a_5547_975.t5 a_5547_975.t3 285.986
R20618 a_5547_975.n0 a_5547_975.t4 282.573
R20619 a_5547_975.n1 a_5547_975.t0 202.857
R20620 a_5547_975.n1 a_5547_975.n0 173.817
R20621 a_5547_975.n1 a_5547_975.t1 20.826
R20622 a_5547_975.n2 a_5547_975.n1 20.689
R20623 a_3152_678.n0 a_3152_678.t2 362.857
R20624 a_3152_678.t3 a_3152_678.t5 337.399
R20625 a_3152_678.t5 a_3152_678.t4 298.839
R20626 a_3152_678.n0 a_3152_678.t3 280.405
R20627 a_3152_678.n1 a_3152_678.t0 200
R20628 a_3152_678.n1 a_3152_678.n0 172.311
R20629 a_3152_678.n2 a_3152_678.n1 24
R20630 a_3152_678.n1 a_3152_678.t1 21.212
R20631 a_8221_n5850.n0 a_8221_n5850.t4 1465.51
R20632 a_8221_n5850.n0 a_8221_n5850.t3 712.44
R20633 a_8221_n5850.n1 a_8221_n5850.t0 375.067
R20634 a_8221_n5850.n1 a_8221_n5850.t1 272.668
R20635 a_8221_n5850.n2 a_8221_n5850.n0 143.764
R20636 a_8221_n5850.t2 a_8221_n5850.n2 78.193
R20637 a_8221_n5850.n2 a_8221_n5850.n1 4.517
R20638 a_1522_4148.n0 a_1522_4148.t1 358.166
R20639 a_1522_4148.t3 a_1522_4148.t5 337.399
R20640 a_1522_4148.t5 a_1522_4148.t4 285.986
R20641 a_1522_4148.n0 a_1522_4148.t3 282.573
R20642 a_1522_4148.n1 a_1522_4148.t2 202.857
R20643 a_1522_4148.n1 a_1522_4148.n0 173.817
R20644 a_1522_4148.n1 a_1522_4148.t0 20.826
R20645 a_1522_4148.n2 a_1522_4148.n1 20.689
R20646 a_8997_2943.n0 a_8997_2943.t2 358.166
R20647 a_8997_2943.t4 a_8997_2943.t5 337.399
R20648 a_8997_2943.t5 a_8997_2943.t3 285.986
R20649 a_8997_2943.n0 a_8997_2943.t4 282.573
R20650 a_8997_2943.n1 a_8997_2943.t0 202.857
R20651 a_8997_2943.n1 a_8997_2943.n0 173.817
R20652 a_8997_2943.n1 a_8997_2943.t1 20.826
R20653 a_8997_2943.n2 a_8997_2943.n1 20.689
R20654 a_3617_1698.t0 a_3617_1698.t1 242.857
R20655 a_6697_n30.n0 a_6697_n30.t1 358.166
R20656 a_6697_n30.t5 a_6697_n30.t3 337.399
R20657 a_6697_n30.t3 a_6697_n30.t4 285.986
R20658 a_6697_n30.n0 a_6697_n30.t5 282.573
R20659 a_6697_n30.n1 a_6697_n30.t0 202.857
R20660 a_6697_n30.n1 a_6697_n30.n0 173.817
R20661 a_6697_n30.n1 a_6697_n30.t2 20.826
R20662 a_6697_n30.n2 a_6697_n30.n1 20.689
R20663 a_6602_n45.n0 a_6602_n45.t1 362.857
R20664 a_6602_n45.t3 a_6602_n45.t5 337.399
R20665 a_6602_n45.t5 a_6602_n45.t4 298.839
R20666 a_6602_n45.n0 a_6602_n45.t3 280.405
R20667 a_6602_n45.n1 a_6602_n45.t2 200
R20668 a_6602_n45.n1 a_6602_n45.n0 172.311
R20669 a_6602_n45.n2 a_6602_n45.n1 24
R20670 a_6602_n45.n1 a_6602_n45.t0 21.212
R20671 a_12736_n8026.n0 a_12736_n8026.t0 65.063
R20672 a_12736_n8026.n0 a_12736_n8026.t2 42.011
R20673 a_12736_n8026.t1 a_12736_n8026.n0 2.113
R20674 a_8792_3184.t0 a_8792_3184.t1 242.857
R20675 a_8997_211.n0 a_8997_211.t1 358.166
R20676 a_8997_211.t5 a_8997_211.t4 337.399
R20677 a_8997_211.t4 a_8997_211.t3 285.986
R20678 a_8997_211.n0 a_8997_211.t5 282.573
R20679 a_8997_211.n1 a_8997_211.t2 202.857
R20680 a_8997_211.n1 a_8997_211.n0 173.817
R20681 a_8997_211.n1 a_8997_211.t0 20.826
R20682 a_8997_211.n2 a_8997_211.n1 20.689
R20683 a_9405_n8583.n0 a_9405_n8583.t4 1465.51
R20684 a_9405_n8583.n0 a_9405_n8583.t3 712.44
R20685 a_9405_n8583.n1 a_9405_n8583.t0 375.067
R20686 a_9405_n8583.n1 a_9405_n8583.t1 272.668
R20687 a_9405_n8583.n2 a_9405_n8583.n0 143.764
R20688 a_9405_n8583.t2 a_9405_n8583.n2 78.193
R20689 a_9405_n8583.n2 a_9405_n8583.n1 4.517
R20690 a_6602_2406.n0 a_6602_2406.t0 362.857
R20691 a_6602_2406.t3 a_6602_2406.t5 337.399
R20692 a_6602_2406.t5 a_6602_2406.t4 298.839
R20693 a_6602_2406.n0 a_6602_2406.t3 280.405
R20694 a_6602_2406.n1 a_6602_2406.t2 200
R20695 a_6602_2406.n1 a_6602_2406.n0 172.311
R20696 a_6602_2406.n2 a_6602_2406.n1 24
R20697 a_6602_2406.n1 a_6602_2406.t1 21.212
R20698 a_8422_693.n0 a_8422_693.t1 358.166
R20699 a_8422_693.t3 a_8422_693.t5 337.399
R20700 a_8422_693.t5 a_8422_693.t4 285.986
R20701 a_8422_693.n0 a_8422_693.t3 282.573
R20702 a_8422_693.n1 a_8422_693.t2 202.857
R20703 a_8422_693.n1 a_8422_693.n0 173.817
R20704 a_8422_693.n1 a_8422_693.t0 20.826
R20705 a_8422_693.n2 a_8422_693.n1 20.689
R20706 a_4675_n8583.n0 a_4675_n8583.t3 1465.51
R20707 a_4675_n8583.n0 a_4675_n8583.t4 712.44
R20708 a_4675_n8583.n1 a_4675_n8583.t0 375.067
R20709 a_4675_n8583.n1 a_4675_n8583.t2 272.668
R20710 a_4675_n8583.n2 a_4675_n8583.n0 143.764
R20711 a_4675_n8583.t1 a_4675_n8583.n2 78.193
R20712 a_4675_n8583.n2 a_4675_n8583.n1 4.517
R20713 a_8902_3410.n0 a_8902_3410.t1 362.857
R20714 a_8902_3410.t5 a_8902_3410.t4 337.399
R20715 a_8902_3410.t4 a_8902_3410.t3 298.839
R20716 a_8902_3410.n0 a_8902_3410.t5 280.405
R20717 a_8902_3410.n1 a_8902_3410.t0 200
R20718 a_8902_3410.n1 a_8902_3410.n0 172.311
R20719 a_8902_3410.n2 a_8902_3410.n1 24
R20720 a_8902_3410.n1 a_8902_3410.t2 21.212
R20721 a_8915_3425.t0 a_8915_3425.t1 242.857
R20722 a_2672_2421.n0 a_2672_2421.t0 358.166
R20723 a_2672_2421.t3 a_2672_2421.t4 337.399
R20724 a_2672_2421.t4 a_2672_2421.t5 285.986
R20725 a_2672_2421.n0 a_2672_2421.t3 282.573
R20726 a_2672_2421.n1 a_2672_2421.t2 202.857
R20727 a_2672_2421.n1 a_2672_2421.n0 173.817
R20728 a_2672_2421.n1 a_2672_2421.t1 20.826
R20729 a_2672_2421.n2 a_2672_2421.n1 20.689
R20730 a_2577_2406.n0 a_2577_2406.t1 362.857
R20731 a_2577_2406.t3 a_2577_2406.t4 337.399
R20732 a_2577_2406.t4 a_2577_2406.t5 298.839
R20733 a_2577_2406.n0 a_2577_2406.t3 280.405
R20734 a_2577_2406.n1 a_2577_2406.t2 200
R20735 a_2577_2406.n1 a_2577_2406.n0 172.311
R20736 a_2577_2406.n2 a_2577_2406.n1 24
R20737 a_2577_2406.n1 a_2577_2406.t0 21.212
R20738 a_6040_975.t0 a_6040_975.t1 242.857
R20739 a_7067_n30.t0 a_7067_n30.t1 242.857
R20740 a_4972_2943.n0 a_4972_2943.t2 358.166
R20741 a_4972_2943.t3 a_4972_2943.t5 337.399
R20742 a_4972_2943.t5 a_4972_2943.t4 285.986
R20743 a_4972_2943.n0 a_4972_2943.t3 282.573
R20744 a_4972_2943.n1 a_4972_2943.t0 202.857
R20745 a_4972_2943.n1 a_4972_2943.n0 173.817
R20746 a_4972_2943.n1 a_4972_2943.t1 20.826
R20747 a_4972_2943.n2 a_4972_2943.n1 20.689
R20748 a_4877_2928.n0 a_4877_2928.t2 362.857
R20749 a_4877_2928.t4 a_4877_2928.t3 337.399
R20750 a_4877_2928.t3 a_4877_2928.t5 298.839
R20751 a_4877_2928.n0 a_4877_2928.t4 280.405
R20752 a_4877_2928.n1 a_4877_2928.t0 200
R20753 a_4877_2928.n1 a_4877_2928.n0 172.311
R20754 a_4877_2928.n2 a_4877_2928.n1 24
R20755 a_4877_2928.n1 a_4877_2928.t1 21.212
R20756 RWL[7].n0 RWL[7].t10 154.243
R20757 RWL[7].n14 RWL[7].t0 149.249
R20758 RWL[7].n13 RWL[7].t5 149.249
R20759 RWL[7].n12 RWL[7].t12 149.249
R20760 RWL[7].n11 RWL[7].t1 149.249
R20761 RWL[7].n10 RWL[7].t14 149.249
R20762 RWL[7].n9 RWL[7].t6 149.249
R20763 RWL[7].n8 RWL[7].t13 149.249
R20764 RWL[7].n7 RWL[7].t3 149.249
R20765 RWL[7].n6 RWL[7].t15 149.249
R20766 RWL[7].n5 RWL[7].t9 149.249
R20767 RWL[7].n4 RWL[7].t2 149.249
R20768 RWL[7].n3 RWL[7].t7 149.249
R20769 RWL[7].n2 RWL[7].t8 149.249
R20770 RWL[7].n1 RWL[7].t11 149.249
R20771 RWL[7].n0 RWL[7].t4 149.249
R20772 RWL[7] RWL[7].n14 42.872
R20773 RWL[7].n1 RWL[7].n0 4.994
R20774 RWL[7].n2 RWL[7].n1 4.994
R20775 RWL[7].n3 RWL[7].n2 4.994
R20776 RWL[7].n4 RWL[7].n3 4.994
R20777 RWL[7].n5 RWL[7].n4 4.994
R20778 RWL[7].n6 RWL[7].n5 4.994
R20779 RWL[7].n7 RWL[7].n6 4.994
R20780 RWL[7].n8 RWL[7].n7 4.994
R20781 RWL[7].n9 RWL[7].n8 4.994
R20782 RWL[7].n10 RWL[7].n9 4.994
R20783 RWL[7].n11 RWL[7].n10 4.994
R20784 RWL[7].n12 RWL[7].n11 4.994
R20785 RWL[7].n13 RWL[7].n12 4.994
R20786 RWL[7].n14 RWL[7].n13 4.994
R20787 a_290_1939.t0 a_290_1939.t1 242.857
R20788 a_7752_2165.n0 a_7752_2165.t2 362.857
R20789 a_7752_2165.t3 a_7752_2165.t4 337.399
R20790 a_7752_2165.t4 a_7752_2165.t5 298.839
R20791 a_7752_2165.n0 a_7752_2165.t3 280.405
R20792 a_7752_2165.n1 a_7752_2165.t0 200
R20793 a_7752_2165.n1 a_7752_2165.n0 172.311
R20794 a_7752_2165.n2 a_7752_2165.n1 24
R20795 a_7752_2165.n1 a_7752_2165.t1 21.212
R20796 a_9367_2943.t0 a_9367_2943.t1 242.857
R20797 a_4192_1939.t0 a_4192_1939.t1 242.857
R20798 a_3740_3907.t0 a_3740_3907.t1 242.857
R20799 a_4745_n8071.n0 a_4745_n8071.t0 63.08
R20800 a_4745_n8071.n0 a_4745_n8071.t2 41.307
R20801 a_4745_n8071.t1 a_4745_n8071.n0 2.251
R20802 RWL[11].n0 RWL[11].t14 154.243
R20803 RWL[11].n14 RWL[11].t4 149.249
R20804 RWL[11].n13 RWL[11].t9 149.249
R20805 RWL[11].n12 RWL[11].t0 149.249
R20806 RWL[11].n11 RWL[11].t5 149.249
R20807 RWL[11].n10 RWL[11].t2 149.249
R20808 RWL[11].n9 RWL[11].t10 149.249
R20809 RWL[11].n8 RWL[11].t1 149.249
R20810 RWL[11].n7 RWL[11].t7 149.249
R20811 RWL[11].n6 RWL[11].t3 149.249
R20812 RWL[11].n5 RWL[11].t13 149.249
R20813 RWL[11].n4 RWL[11].t6 149.249
R20814 RWL[11].n3 RWL[11].t11 149.249
R20815 RWL[11].n2 RWL[11].t12 149.249
R20816 RWL[11].n1 RWL[11].t15 149.249
R20817 RWL[11].n0 RWL[11].t8 149.249
R20818 RWL[11] RWL[11].n14 42.872
R20819 RWL[11].n1 RWL[11].n0 4.994
R20820 RWL[11].n2 RWL[11].n1 4.994
R20821 RWL[11].n3 RWL[11].n2 4.994
R20822 RWL[11].n4 RWL[11].n3 4.994
R20823 RWL[11].n5 RWL[11].n4 4.994
R20824 RWL[11].n6 RWL[11].n5 4.994
R20825 RWL[11].n7 RWL[11].n6 4.994
R20826 RWL[11].n8 RWL[11].n7 4.994
R20827 RWL[11].n9 RWL[11].n8 4.994
R20828 RWL[11].n10 RWL[11].n9 4.994
R20829 RWL[11].n11 RWL[11].n10 4.994
R20830 RWL[11].n12 RWL[11].n11 4.994
R20831 RWL[11].n13 RWL[11].n12 4.994
R20832 RWL[11].n14 RWL[11].n13 4.994
R20833 a_1440_975.t0 a_1440_975.t1 242.857
R20834 a_7847_2180.n0 a_7847_2180.t2 358.166
R20835 a_7847_2180.t4 a_7847_2180.t5 337.399
R20836 a_7847_2180.t5 a_7847_2180.t3 285.986
R20837 a_7847_2180.n0 a_7847_2180.t4 282.573
R20838 a_7847_2180.n1 a_7847_2180.t0 202.857
R20839 a_7847_2180.n1 a_7847_2180.n0 173.817
R20840 a_7847_2180.n1 a_7847_2180.t1 20.826
R20841 a_7847_2180.n2 a_7847_2180.n1 20.689
R20842 a_8217_2180.t0 a_8217_2180.t1 242.857
R20843 a_277_1683.n0 a_277_1683.t1 362.857
R20844 a_277_1683.t4 a_277_1683.t5 337.399
R20845 a_277_1683.t5 a_277_1683.t3 298.839
R20846 a_277_1683.n0 a_277_1683.t4 280.405
R20847 a_277_1683.n1 a_277_1683.t2 200
R20848 a_277_1683.n1 a_277_1683.n0 172.311
R20849 a_277_1683.n2 a_277_1683.n1 24
R20850 a_277_1683.n1 a_277_1683.t0 21.212
R20851 a_290_1698.t0 a_290_1698.t1 242.857
R20852 ADC0_OUT[3].n0 ADC0_OUT[3].t3 1355.37
R20853 ADC0_OUT[3].n0 ADC0_OUT[3].t4 820.859
R20854 ADC0_OUT[3].n3 ADC0_OUT[3].t0 342.691
R20855 ADC0_OUT[3].n2 ADC0_OUT[3].t1 266.644
R20856 ADC0_OUT[3].n1 ADC0_OUT[3].n0 149.035
R20857 ADC0_OUT[3].n1 ADC0_OUT[3].t2 45.968
R20858 ADC0_OUT[3].n3 ADC0_OUT[3].n2 41.411
R20859 ADC0_OUT[3] ADC0_OUT[3].n3 22.236
R20860 ADC0_OUT[3].n2 ADC0_OUT[3].n1 17.317
R20861 a_n3495_n8071.n0 a_n3495_n8071.t0 63.08
R20862 a_n3495_n8071.n0 a_n3495_n8071.t2 41.307
R20863 a_n3495_n8071.t1 a_n3495_n8071.n0 2.251
R20864 a_n3565_n8583.n0 a_n3565_n8583.t4 1465.51
R20865 a_n3565_n8583.n0 a_n3565_n8583.t3 712.44
R20866 a_n3565_n8583.n1 a_n3565_n8583.t0 375.067
R20867 a_n3565_n8583.n1 a_n3565_n8583.t2 272.668
R20868 a_n3565_n8583.n2 a_n3565_n8583.n0 143.764
R20869 a_n3565_n8583.t1 a_n3565_n8583.n2 78.193
R20870 a_n3565_n8583.n2 a_n3565_n8583.n1 4.517
R20871 a_4890_n1053.t0 a_4890_n1053.t1 242.857
R20872 a_4192_1698.t0 a_4192_1698.t1 242.857
R20873 a_3042_3666.t0 a_3042_3666.t1 242.857
R20874 a_3617_1216.t0 a_3617_1216.t1 242.857
R20875 a_7109_n8071.n0 a_7109_n8071.t0 63.08
R20876 a_7109_n8071.n0 a_7109_n8071.t2 41.307
R20877 a_7109_n8071.t1 a_7109_n8071.n0 2.251
R20878 SA_OUT[8].n1 SA_OUT[8].t4 661.027
R20879 SA_OUT[8].n1 SA_OUT[8].t3 392.255
R20880 SA_OUT[8].n2 SA_OUT[8].t1 223.716
R20881 SA_OUT[8].n0 SA_OUT[8].t0 153.977
R20882 SA_OUT[8].n2 SA_OUT[8].n1 143.764
R20883 SA_OUT[8].n0 SA_OUT[8].t2 59.86
R20884 SA_OUT[8] SA_OUT[8].n3 15.15
R20885 SA_OUT[8].n3 SA_OUT[8].n0 2.258
R20886 SA_OUT[8].n3 SA_OUT[8].n2 2.258
R20887 a_4910_n1371.n1 a_4910_n1371.t3 550.94
R20888 a_4910_n1371.n1 a_4910_n1371.t4 500.621
R20889 a_4910_n1371.t0 a_4910_n1371.n2 192.787
R20890 a_4910_n1371.n0 a_4910_n1371.t2 163.997
R20891 a_4910_n1371.n2 a_4910_n1371.n1 149.035
R20892 a_4910_n1371.n0 a_4910_n1371.t1 54.068
R20893 a_4910_n1371.n2 a_4910_n1371.n0 17.317
R20894 a_8327_n827.n0 a_8327_n827.t2 362.857
R20895 a_8327_n827.t3 a_8327_n827.t4 337.399
R20896 a_8327_n827.t4 a_8327_n827.t5 298.839
R20897 a_8327_n827.n0 a_8327_n827.t3 280.405
R20898 a_8327_n827.n1 a_8327_n827.t0 200
R20899 a_8327_n827.n1 a_8327_n827.n0 172.311
R20900 a_8327_n827.n2 a_8327_n827.n1 24
R20901 a_8327_n827.n1 a_8327_n827.t1 21.212
R20902 a_4315_3666.t0 a_4315_3666.t1 242.857
R20903 a_5465_1698.t0 a_5465_1698.t1 242.857
R20904 a_8327_1683.n0 a_8327_1683.t2 362.857
R20905 a_8327_1683.t5 a_8327_1683.t3 337.399
R20906 a_8327_1683.t3 a_8327_1683.t4 298.839
R20907 a_8327_1683.n0 a_8327_1683.t5 280.405
R20908 a_8327_1683.n1 a_8327_1683.t0 200
R20909 a_8327_1683.n1 a_8327_1683.n0 172.311
R20910 a_8327_1683.n2 a_8327_1683.n1 24
R20911 a_8327_1683.n1 a_8327_1683.t1 21.212
R20912 a_6777_n7825.t0 a_6777_n7825.t1 42.705
R20913 a_6812_n8026.n0 a_6812_n8026.t0 65.063
R20914 a_6812_n8026.n0 a_6812_n8026.t2 42.011
R20915 a_6812_n8026.t1 a_6812_n8026.n0 2.113
R20916 a_1317_n30.t0 a_1317_n30.t1 242.857
R20917 a_5465_n812.t0 a_5465_n812.t1 242.857
R20918 a_n3792_n3770.n0 a_n3792_n3770.t0 65.064
R20919 a_n3792_n3770.n0 a_n3792_n3770.t2 42.011
R20920 a_n3792_n3770.t1 a_n3792_n3770.n0 2.113
R20921 a_7272_1939.n0 a_7272_1939.t2 358.166
R20922 a_7272_1939.t5 a_7272_1939.t4 337.399
R20923 a_7272_1939.t4 a_7272_1939.t3 285.986
R20924 a_7272_1939.n0 a_7272_1939.t5 282.573
R20925 a_7272_1939.n1 a_7272_1939.t0 202.857
R20926 a_7272_1939.n1 a_7272_1939.n0 173.817
R20927 a_7272_1939.n1 a_7272_1939.t1 20.826
R20928 a_7272_1939.n2 a_7272_1939.n1 20.689
R20929 a_7642_1939.t0 a_7642_1939.t1 242.857
R20930 a_3740_n271.t0 a_3740_n271.t1 242.857
R20931 a_3822_4686.n0 a_3822_4686.t2 358.166
R20932 a_3822_4686.t5 a_3822_4686.t4 337.399
R20933 a_3822_4686.t4 a_3822_4686.t3 285.986
R20934 a_3822_4686.n0 a_3822_4686.t5 282.573
R20935 a_3822_4686.n1 a_3822_4686.t0 202.857
R20936 a_3822_4686.n1 a_3822_4686.n0 173.817
R20937 a_3822_4686.n1 a_3822_4686.t1 20.826
R20938 a_3822_4686.n2 a_3822_4686.n1 20.689
R20939 a_6777_n6849.t0 a_6777_n6849.t1 42.707
R20940 a_7210_n1371.n1 a_7210_n1371.t4 550.94
R20941 a_7210_n1371.n1 a_7210_n1371.t3 500.621
R20942 a_7210_n1371.t1 a_7210_n1371.n2 192.787
R20943 a_7210_n1371.n0 a_7210_n1371.t2 163.997
R20944 a_7210_n1371.n2 a_7210_n1371.n1 149.035
R20945 a_7210_n1371.n0 a_7210_n1371.t0 54.068
R20946 a_7210_n1371.n2 a_7210_n1371.n0 17.317
R20947 a_5465_211.t0 a_5465_211.t1 242.857
R20948 a_3165_n30.t0 a_3165_n30.t1 242.857
R20949 a_n314_n4116.t0 a_n314_n4116.t1 42.707
R20950 a_947_3666.n0 a_947_3666.t0 358.166
R20951 a_947_3666.t5 a_947_3666.t3 337.399
R20952 a_947_3666.t3 a_947_3666.t4 285.986
R20953 a_947_3666.n0 a_947_3666.t5 282.573
R20954 a_947_3666.n1 a_947_3666.t2 202.857
R20955 a_947_3666.n1 a_947_3666.n0 173.817
R20956 a_947_3666.n1 a_947_3666.t1 20.826
R20957 a_947_3666.n2 a_947_3666.n1 20.689
R20958 a_852_3651.n0 a_852_3651.t1 362.857
R20959 a_852_3651.t3 a_852_3651.t4 337.399
R20960 a_852_3651.t4 a_852_3651.t5 298.839
R20961 a_852_3651.n0 a_852_3651.t3 280.405
R20962 a_852_3651.n1 a_852_3651.t2 200
R20963 a_852_3651.n1 a_852_3651.n0 172.311
R20964 a_852_3651.n2 a_852_3651.n1 24
R20965 a_852_3651.n1 a_852_3651.t0 21.212
R20966 a_277_2647.n0 a_277_2647.t1 362.857
R20967 a_277_2647.t3 a_277_2647.t4 337.399
R20968 a_277_2647.t4 a_277_2647.t5 298.839
R20969 a_277_2647.n0 a_277_2647.t3 280.405
R20970 a_277_2647.n1 a_277_2647.t2 200
R20971 a_277_2647.n1 a_277_2647.n0 172.311
R20972 a_277_2647.n2 a_277_2647.n1 24
R20973 a_277_2647.n1 a_277_2647.t0 21.212
R20974 a_7272_2662.n0 a_7272_2662.t0 358.166
R20975 a_7272_2662.t3 a_7272_2662.t5 337.399
R20976 a_7272_2662.t5 a_7272_2662.t4 285.986
R20977 a_7272_2662.n0 a_7272_2662.t3 282.573
R20978 a_7272_2662.n1 a_7272_2662.t2 202.857
R20979 a_7272_2662.n1 a_7272_2662.n0 173.817
R20980 a_7272_2662.n1 a_7272_2662.t1 20.826
R20981 a_7272_2662.n2 a_7272_2662.n1 20.689
R20982 a_7177_2647.n0 a_7177_2647.t1 362.857
R20983 a_7177_2647.t3 a_7177_2647.t4 337.399
R20984 a_7177_2647.t4 a_7177_2647.t5 298.839
R20985 a_7177_2647.n0 a_7177_2647.t3 280.405
R20986 a_7177_2647.n1 a_7177_2647.t2 200
R20987 a_7177_2647.n1 a_7177_2647.n0 172.311
R20988 a_7177_2647.n2 a_7177_2647.n1 24
R20989 a_7177_2647.n1 a_7177_2647.t0 21.212
R20990 a_8915_452.t0 a_8915_452.t1 242.857
R20991 a_7847_2943.n0 a_7847_2943.t2 358.166
R20992 a_7847_2943.t5 a_7847_2943.t3 337.399
R20993 a_7847_2943.t3 a_7847_2943.t4 285.986
R20994 a_7847_2943.n0 a_7847_2943.t5 282.573
R20995 a_7847_2943.n1 a_7847_2943.t0 202.857
R20996 a_7847_2943.n1 a_7847_2943.n0 173.817
R20997 a_7847_2943.n1 a_7847_2943.t1 20.826
R20998 a_7847_2943.n2 a_7847_2943.n1 20.689
R20999 a_2672_1939.n0 a_2672_1939.t2 358.166
R21000 a_2672_1939.t3 a_2672_1939.t4 337.399
R21001 a_2672_1939.t4 a_2672_1939.t5 285.986
R21002 a_2672_1939.n0 a_2672_1939.t3 282.573
R21003 a_2672_1939.n1 a_2672_1939.t0 202.857
R21004 a_2672_1939.n1 a_2672_1939.n0 173.817
R21005 a_2672_1939.n1 a_2672_1939.t1 20.826
R21006 a_2672_1939.n2 a_2672_1939.n1 20.689
R21007 a_947_693.n0 a_947_693.t2 358.166
R21008 a_947_693.t5 a_947_693.t4 337.399
R21009 a_947_693.t4 a_947_693.t3 285.986
R21010 a_947_693.n0 a_947_693.t5 282.573
R21011 a_947_693.n1 a_947_693.t0 202.857
R21012 a_947_693.n1 a_947_693.n0 173.817
R21013 a_947_693.n1 a_947_693.t1 20.826
R21014 a_947_693.n2 a_947_693.n1 20.689
R21015 a_8291_n5338.n0 a_8291_n5338.t0 63.08
R21016 a_8291_n5338.n0 a_8291_n5338.t2 41.307
R21017 a_8291_n5338.t1 a_8291_n5338.n0 2.251
R21018 a_8291_n4470.n0 a_8291_n4470.t0 63.08
R21019 a_8291_n4470.n0 a_8291_n4470.t2 41.305
R21020 a_8291_n4470.t1 a_8291_n4470.n0 2.251
R21021 a_3740_3425.t0 a_3740_3425.t1 242.857
R21022 a_4890_1457.t0 a_4890_1457.t1 242.857
R21023 a_372_1939.n0 a_372_1939.t1 358.166
R21024 a_372_1939.t4 a_372_1939.t3 337.399
R21025 a_372_1939.t3 a_372_1939.t5 285.986
R21026 a_372_1939.n0 a_372_1939.t4 282.573
R21027 a_372_1939.n1 a_372_1939.t2 202.857
R21028 a_372_1939.n1 a_372_1939.n0 173.817
R21029 a_372_1939.n1 a_372_1939.t0 20.826
R21030 a_372_1939.n2 a_372_1939.n1 20.689
R21031 a_277_1924.n0 a_277_1924.t1 362.857
R21032 a_277_1924.t5 a_277_1924.t3 337.399
R21033 a_277_1924.t3 a_277_1924.t4 298.839
R21034 a_277_1924.n0 a_277_1924.t5 280.405
R21035 a_277_1924.n1 a_277_1924.t2 200
R21036 a_277_1924.n1 a_277_1924.n0 172.311
R21037 a_277_1924.n2 a_277_1924.n1 24
R21038 a_277_1924.n1 a_277_1924.t0 21.212
R21039 a_2097_n812.n0 a_2097_n812.t1 358.166
R21040 a_2097_n812.t5 a_2097_n812.t3 337.399
R21041 a_2097_n812.t3 a_2097_n812.t4 285.986
R21042 a_2097_n812.n0 a_2097_n812.t5 282.573
R21043 a_2097_n812.n1 a_2097_n812.t0 202.857
R21044 a_2097_n812.n1 a_2097_n812.n0 173.817
R21045 a_2097_n812.n1 a_2097_n812.t2 20.826
R21046 a_2097_n812.n2 a_2097_n812.n1 20.689
R21047 a_2002_n827.n0 a_2002_n827.t2 362.857
R21048 a_2002_n827.t3 a_2002_n827.t5 337.399
R21049 a_2002_n827.t5 a_2002_n827.t4 298.839
R21050 a_2002_n827.n0 a_2002_n827.t3 280.405
R21051 a_2002_n827.n1 a_2002_n827.t0 200
R21052 a_2002_n827.n1 a_2002_n827.n0 172.311
R21053 a_2002_n827.n2 a_2002_n827.n1 24
R21054 a_2002_n827.n1 a_2002_n827.t1 21.212
R21055 a_7642_1698.t0 a_7642_1698.t1 242.857
R21056 a_6602_437.n0 a_6602_437.t2 362.857
R21057 a_6602_437.t4 a_6602_437.t3 337.399
R21058 a_6602_437.t3 a_6602_437.t5 298.839
R21059 a_6602_437.n0 a_6602_437.t4 280.405
R21060 a_6602_437.n1 a_6602_437.t0 200
R21061 a_6602_437.n1 a_6602_437.n0 172.311
R21062 a_6602_437.n2 a_6602_437.n1 24
R21063 a_6602_437.n1 a_6602_437.t1 21.212
R21064 a_290_1216.t0 a_290_1216.t1 242.857
R21065 a_1427_1683.n0 a_1427_1683.t1 362.857
R21066 a_1427_1683.t3 a_1427_1683.t4 337.399
R21067 a_1427_1683.t4 a_1427_1683.t5 298.839
R21068 a_1427_1683.n0 a_1427_1683.t3 280.405
R21069 a_1427_1683.n1 a_1427_1683.t0 200
R21070 a_1427_1683.n1 a_1427_1683.n0 172.311
R21071 a_1427_1683.n2 a_1427_1683.n1 24
R21072 a_1427_1683.n1 a_1427_1683.t2 21.212
R21073 a_2311_n4483.n0 a_2311_n4483.t3 1464.36
R21074 a_2311_n4483.n0 a_2311_n4483.t4 713.588
R21075 a_2311_n4483.n1 a_2311_n4483.t0 374.998
R21076 a_2311_n4483.n1 a_2311_n4483.t2 273.351
R21077 a_2311_n4483.n2 a_2311_n4483.n0 143.764
R21078 a_2311_n4483.t1 a_2311_n4483.n2 78.209
R21079 a_2311_n4483.n2 a_2311_n4483.n1 4.517
R21080 a_372_2662.n0 a_372_2662.t1 358.166
R21081 a_372_2662.t5 a_372_2662.t4 337.399
R21082 a_372_2662.t4 a_372_2662.t3 285.986
R21083 a_372_2662.n0 a_372_2662.t5 282.573
R21084 a_372_2662.n1 a_372_2662.t2 202.857
R21085 a_372_2662.n1 a_372_2662.n0 173.817
R21086 a_372_2662.n1 a_372_2662.t0 20.826
R21087 a_372_2662.n2 a_372_2662.n1 20.689
R21088 a_742_2662.t0 a_742_2662.t1 242.857
R21089 a_8915_1698.t0 a_8915_1698.t1 242.857
R21090 a_4192_1216.t0 a_4192_1216.t1 242.857
R21091 a_4397_211.n0 a_4397_211.t2 358.166
R21092 a_4397_211.t5 a_4397_211.t4 337.399
R21093 a_4397_211.t4 a_4397_211.t3 285.986
R21094 a_4397_211.n0 a_4397_211.t5 282.573
R21095 a_4397_211.n1 a_4397_211.t0 202.857
R21096 a_4397_211.n1 a_4397_211.n0 173.817
R21097 a_4397_211.n1 a_4397_211.t1 20.826
R21098 a_4397_211.n2 a_4397_211.n1 20.689
R21099 SA_OUT[9].n0 SA_OUT[9].t3 661.027
R21100 SA_OUT[9].n0 SA_OUT[9].t4 392.255
R21101 SA_OUT[9].n1 SA_OUT[9].t1 223.716
R21102 SA_OUT[9].n2 SA_OUT[9].t2 153.977
R21103 SA_OUT[9].n1 SA_OUT[9].n0 143.764
R21104 SA_OUT[9].n2 SA_OUT[9].t0 59.86
R21105 SA_OUT[9] SA_OUT[9].n2 14.841
R21106 SA_OUT[9].n2 SA_OUT[9].n1 4.517
R21107 a_5485_n1371.n1 a_5485_n1371.t4 550.94
R21108 a_5485_n1371.n1 a_5485_n1371.t3 500.621
R21109 a_5485_n1371.t1 a_5485_n1371.n2 192.787
R21110 a_5485_n1371.n0 a_5485_n1371.t0 163.997
R21111 a_5485_n1371.n2 a_5485_n1371.n1 149.035
R21112 a_5485_n1371.n0 a_5485_n1371.t2 54.068
R21113 a_5485_n1371.n2 a_5485_n1371.n0 17.317
R21114 a_5577_n1770.t0 a_5577_n1770.n0 182.779
R21115 a_5577_n1770.n0 a_5577_n1770.t1 111.474
R21116 a_7765_n1053.t0 a_7765_n1053.t1 242.857
R21117 ADC11_OUT[0].n0 ADC11_OUT[0].t4 1354.27
R21118 ADC11_OUT[0].n0 ADC11_OUT[0].t3 821.954
R21119 ADC11_OUT[0].n3 ADC11_OUT[0].t0 347.891
R21120 ADC11_OUT[0].n2 ADC11_OUT[0].t2 266.575
R21121 ADC11_OUT[0].n1 ADC11_OUT[0].n0 149.035
R21122 ADC11_OUT[0] ADC11_OUT[0].n3 61.793
R21123 ADC11_OUT[0].n1 ADC11_OUT[0].t1 46.723
R21124 ADC11_OUT[0].n3 ADC11_OUT[0].n2 36.141
R21125 ADC11_OUT[0].n2 ADC11_OUT[0].n1 17.317
R21126 a_9405_n4483.n0 a_9405_n4483.t3 1464.36
R21127 a_9405_n4483.n0 a_9405_n4483.t4 713.588
R21128 a_9405_n4483.n1 a_9405_n4483.t0 374.998
R21129 a_9405_n4483.n1 a_9405_n4483.t1 273.351
R21130 a_9405_n4483.n2 a_9405_n4483.n0 143.764
R21131 a_9405_n4483.t2 a_9405_n4483.n2 78.209
R21132 a_9405_n4483.n2 a_9405_n4483.n1 4.517
R21133 a_6060_n1371.n1 a_6060_n1371.t3 550.94
R21134 a_6060_n1371.n1 a_6060_n1371.t4 500.621
R21135 a_6060_n1371.t1 a_6060_n1371.n2 192.787
R21136 a_6060_n1371.n0 a_6060_n1371.t0 163.997
R21137 a_6060_n1371.n2 a_6060_n1371.n1 149.035
R21138 a_6060_n1371.n0 a_6060_n1371.t2 54.068
R21139 a_6060_n1371.n2 a_6060_n1371.n0 17.317
R21140 a_5465_1216.t0 a_5465_1216.t1 242.857
R21141 a_8327_1201.n0 a_8327_1201.t2 362.857
R21142 a_8327_1201.t5 a_8327_1201.t3 337.399
R21143 a_8327_1201.t3 a_8327_1201.t4 298.839
R21144 a_8327_1201.n0 a_8327_1201.t5 280.405
R21145 a_8327_1201.n1 a_8327_1201.t0 200
R21146 a_8327_1201.n1 a_8327_1201.n0 172.311
R21147 a_8327_1201.n2 a_8327_1201.n1 24
R21148 a_8327_1201.n1 a_8327_1201.t1 21.212
R21149 a_3042_n30.t0 a_3042_n30.t1 242.857
R21150 a_8915_n812.t0 a_8915_n812.t1 242.857
R21151 a_6697_2421.n0 a_6697_2421.t2 358.166
R21152 a_6697_2421.t3 a_6697_2421.t4 337.399
R21153 a_6697_2421.t4 a_6697_2421.t5 285.986
R21154 a_6697_2421.n0 a_6697_2421.t3 282.573
R21155 a_6697_2421.n1 a_6697_2421.t0 202.857
R21156 a_6697_2421.n1 a_6697_2421.n0 173.817
R21157 a_6697_2421.n1 a_6697_2421.t1 20.826
R21158 a_6697_2421.n2 a_6697_2421.n1 20.689
R21159 a_8488_n6847.t1 a_8488_n6847.t0 336.812
R21160 a_8429_n7203.t0 a_8429_n7203.t1 68.741
R21161 RWLB[9].n0 RWLB[9].t3 154.228
R21162 RWLB[9].n14 RWLB[9].t4 149.249
R21163 RWLB[9].n13 RWLB[9].t6 149.249
R21164 RWLB[9].n12 RWLB[9].t1 149.249
R21165 RWLB[9].n11 RWLB[9].t11 149.249
R21166 RWLB[9].n10 RWLB[9].t5 149.249
R21167 RWLB[9].n9 RWLB[9].t8 149.249
R21168 RWLB[9].n8 RWLB[9].t9 149.249
R21169 RWLB[9].n7 RWLB[9].t14 149.249
R21170 RWLB[9].n6 RWLB[9].t7 149.249
R21171 RWLB[9].n5 RWLB[9].t12 149.249
R21172 RWLB[9].n4 RWLB[9].t13 149.249
R21173 RWLB[9].n3 RWLB[9].t2 149.249
R21174 RWLB[9].n2 RWLB[9].t10 149.249
R21175 RWLB[9].n1 RWLB[9].t0 149.249
R21176 RWLB[9].n0 RWLB[9].t15 149.249
R21177 RWLB[9] RWLB[9].n14 47.816
R21178 RWLB[9].n1 RWLB[9].n0 4.979
R21179 RWLB[9].n2 RWLB[9].n1 4.979
R21180 RWLB[9].n3 RWLB[9].n2 4.979
R21181 RWLB[9].n4 RWLB[9].n3 4.979
R21182 RWLB[9].n5 RWLB[9].n4 4.979
R21183 RWLB[9].n6 RWLB[9].n5 4.979
R21184 RWLB[9].n7 RWLB[9].n6 4.979
R21185 RWLB[9].n8 RWLB[9].n7 4.979
R21186 RWLB[9].n9 RWLB[9].n8 4.979
R21187 RWLB[9].n10 RWLB[9].n9 4.979
R21188 RWLB[9].n11 RWLB[9].n10 4.979
R21189 RWLB[9].n12 RWLB[9].n11 4.979
R21190 RWLB[9].n13 RWLB[9].n12 4.979
R21191 RWLB[9].n14 RWLB[9].n13 4.979
R21192 a_8217_1457.t0 a_8217_1457.t1 242.857
R21193 a_7190_452.t0 a_7190_452.t1 242.857
R21194 a_2002_1924.n0 a_2002_1924.t1 362.857
R21195 a_2002_1924.t3 a_2002_1924.t5 337.399
R21196 a_2002_1924.t5 a_2002_1924.t4 298.839
R21197 a_2002_1924.n0 a_2002_1924.t3 280.405
R21198 a_2002_1924.n1 a_2002_1924.t0 200
R21199 a_2002_1924.n1 a_2002_1924.n0 172.311
R21200 a_2002_1924.n2 a_2002_1924.n1 24
R21201 a_2002_1924.n1 a_2002_1924.t2 21.212
R21202 a_5547_1698.n0 a_5547_1698.t0 358.166
R21203 a_5547_1698.t5 a_5547_1698.t3 337.399
R21204 a_5547_1698.t3 a_5547_1698.t4 285.986
R21205 a_5547_1698.n0 a_5547_1698.t5 282.573
R21206 a_5547_1698.n1 a_5547_1698.t2 202.857
R21207 a_5547_1698.n1 a_5547_1698.n0 173.817
R21208 a_5547_1698.n1 a_5547_1698.t1 20.826
R21209 a_5547_1698.n2 a_5547_1698.n1 20.689
R21210 a_5452_1683.n0 a_5452_1683.t2 362.857
R21211 a_5452_1683.t3 a_5452_1683.t4 337.399
R21212 a_5452_1683.t4 a_5452_1683.t5 298.839
R21213 a_5452_1683.n0 a_5452_1683.t3 280.405
R21214 a_5452_1683.n1 a_5452_1683.t0 200
R21215 a_5452_1683.n1 a_5452_1683.n0 172.311
R21216 a_5452_1683.n2 a_5452_1683.n1 24
R21217 a_5452_1683.n1 a_5452_1683.t1 21.212
R21218 a_3727_2928.n0 a_3727_2928.t2 362.857
R21219 a_3727_2928.t5 a_3727_2928.t3 337.399
R21220 a_3727_2928.t3 a_3727_2928.t4 298.839
R21221 a_3727_2928.n0 a_3727_2928.t5 280.405
R21222 a_3727_2928.n1 a_3727_2928.t0 200
R21223 a_3727_2928.n1 a_3727_2928.n0 172.311
R21224 a_3727_2928.n2 a_3727_2928.n1 24
R21225 a_3727_2928.n1 a_3727_2928.t1 21.212
R21226 SA_OUT[14].n1 SA_OUT[14].t3 661.027
R21227 SA_OUT[14].n1 SA_OUT[14].t4 392.255
R21228 SA_OUT[14].n2 SA_OUT[14].t2 223.716
R21229 SA_OUT[14].n0 SA_OUT[14].t0 153.977
R21230 SA_OUT[14].n2 SA_OUT[14].n1 143.764
R21231 SA_OUT[14].n0 SA_OUT[14].t1 59.86
R21232 SA_OUT[14] SA_OUT[14].n3 13.455
R21233 SA_OUT[14].n3 SA_OUT[14].n2 3.764
R21234 SA_OUT[14].n3 SA_OUT[14].n0 0.752
R21235 a_8360_n1371.n1 a_8360_n1371.t4 550.94
R21236 a_8360_n1371.n1 a_8360_n1371.t3 500.621
R21237 a_8360_n1371.t0 a_8360_n1371.n2 192.787
R21238 a_8360_n1371.n0 a_8360_n1371.t2 163.997
R21239 a_8360_n1371.n2 a_8360_n1371.n1 149.035
R21240 a_8360_n1371.n0 a_8360_n1371.t1 54.068
R21241 a_8360_n1371.n2 a_8360_n1371.n0 17.317
R21242 a_4335_n1371.n1 a_4335_n1371.t3 550.94
R21243 a_4335_n1371.n1 a_4335_n1371.t4 500.621
R21244 a_4335_n1371.t0 a_4335_n1371.n2 192.787
R21245 a_4335_n1371.n0 a_4335_n1371.t2 163.997
R21246 a_4335_n1371.n2 a_4335_n1371.n1 149.035
R21247 a_4335_n1371.n0 a_4335_n1371.t1 54.068
R21248 a_4335_n1371.n2 a_4335_n1371.n0 17.317
R21249 a_5547_n812.n0 a_5547_n812.t1 358.166
R21250 a_5547_n812.t5 a_5547_n812.t3 337.399
R21251 a_5547_n812.t3 a_5547_n812.t4 285.986
R21252 a_5547_n812.n0 a_5547_n812.t5 282.573
R21253 a_5547_n812.n1 a_5547_n812.t0 202.857
R21254 a_5547_n812.n1 a_5547_n812.n0 173.817
R21255 a_5547_n812.n1 a_5547_n812.t2 20.826
R21256 a_5547_n812.n2 a_5547_n812.n1 20.689
R21257 a_5452_n827.n0 a_5452_n827.t2 362.857
R21258 a_5452_n827.t3 a_5452_n827.t4 337.399
R21259 a_5452_n827.t4 a_5452_n827.t5 298.839
R21260 a_5452_n827.n0 a_5452_n827.t3 280.405
R21261 a_5452_n827.n1 a_5452_n827.t0 200
R21262 a_5452_n827.n1 a_5452_n827.n0 172.311
R21263 a_5452_n827.n2 a_5452_n827.n1 24
R21264 a_5452_n827.n1 a_5452_n827.t1 21.212
R21265 a_3617_4445.t0 a_3617_4445.t1 242.857
R21266 a_372_2180.n0 a_372_2180.t0 358.166
R21267 a_372_2180.t3 a_372_2180.t5 337.399
R21268 a_372_2180.t5 a_372_2180.t4 285.986
R21269 a_372_2180.n0 a_372_2180.t3 282.573
R21270 a_372_2180.n1 a_372_2180.t2 202.857
R21271 a_372_2180.n1 a_372_2180.n0 173.817
R21272 a_372_2180.n1 a_372_2180.t1 20.826
R21273 a_372_2180.n2 a_372_2180.n1 20.689
R21274 a_277_2165.n0 a_277_2165.t2 362.857
R21275 a_277_2165.t3 a_277_2165.t4 337.399
R21276 a_277_2165.t4 a_277_2165.t5 298.839
R21277 a_277_2165.n0 a_277_2165.t3 280.405
R21278 a_277_2165.n1 a_277_2165.t0 200
R21279 a_277_2165.n1 a_277_2165.n0 172.311
R21280 a_277_2165.n2 a_277_2165.n1 24
R21281 a_277_2165.n1 a_277_2165.t1 21.212
R21282 a_7642_1216.t0 a_7642_1216.t1 242.857
R21283 a_4302_3651.n0 a_4302_3651.t0 362.857
R21284 a_4302_3651.t3 a_4302_3651.t5 337.399
R21285 a_4302_3651.t5 a_4302_3651.t4 298.839
R21286 a_4302_3651.n0 a_4302_3651.t3 280.405
R21287 a_4302_3651.n1 a_4302_3651.t2 200
R21288 a_4302_3651.n1 a_4302_3651.n0 172.311
R21289 a_4302_3651.n2 a_4302_3651.n1 24
R21290 a_4302_3651.n1 a_4302_3651.t1 21.212
R21291 a_12963_n4483.n0 a_12963_n4483.t4 1464.36
R21292 a_12963_n4483.n0 a_12963_n4483.t3 713.588
R21293 a_12963_n4483.n1 a_12963_n4483.t0 374.998
R21294 a_12963_n4483.n1 a_12963_n4483.t2 273.351
R21295 a_12963_n4483.n2 a_12963_n4483.n0 143.764
R21296 a_12963_n4483.t1 a_12963_n4483.n2 78.209
R21297 a_12963_n4483.n2 a_12963_n4483.n1 4.517
R21298 ADC14_OUT[0].n0 ADC14_OUT[0].t3 1354.27
R21299 ADC14_OUT[0].n0 ADC14_OUT[0].t4 821.954
R21300 ADC14_OUT[0].n3 ADC14_OUT[0].t0 350.15
R21301 ADC14_OUT[0].n2 ADC14_OUT[0].t2 266.575
R21302 ADC14_OUT[0].n1 ADC14_OUT[0].n0 149.035
R21303 ADC14_OUT[0] ADC14_OUT[0].n3 61.534
R21304 ADC14_OUT[0].n1 ADC14_OUT[0].t1 46.723
R21305 ADC14_OUT[0].n3 ADC14_OUT[0].n2 33.882
R21306 ADC14_OUT[0].n2 ADC14_OUT[0].n1 17.317
R21307 a_3042_n1053.t0 a_3042_n1053.t1 242.857
R21308 a_7765_n512.t0 a_7765_n512.t1 242.857
R21309 a_1427_1201.n0 a_1427_1201.t1 362.857
R21310 a_1427_1201.t3 a_1427_1201.t4 337.399
R21311 a_1427_1201.t4 a_1427_1201.t5 298.839
R21312 a_1427_1201.n0 a_1427_1201.t3 280.405
R21313 a_1427_1201.n1 a_1427_1201.t0 200
R21314 a_1427_1201.n1 a_1427_1201.n0 172.311
R21315 a_1427_1201.n2 a_1427_1201.n1 24
R21316 a_1427_1201.n1 a_1427_1201.t2 21.212
R21317 a_453_n2086.t0 a_453_n2086.t1 34.8
R21318 a_8340_3666.t0 a_8340_3666.t1 242.857
R21319 a_8915_1216.t0 a_8915_1216.t1 242.857
R21320 a_7067_452.t0 a_7067_452.t1 242.857
R21321 a_3247_n30.n0 a_3247_n30.t2 358.166
R21322 a_3247_n30.t4 a_3247_n30.t3 337.399
R21323 a_3247_n30.t3 a_3247_n30.t5 285.986
R21324 a_3247_n30.n0 a_3247_n30.t4 282.573
R21325 a_3247_n30.n1 a_3247_n30.t0 202.857
R21326 a_3247_n30.n1 a_3247_n30.n0 173.817
R21327 a_3247_n30.n1 a_3247_n30.t1 20.826
R21328 a_3247_n30.n2 a_3247_n30.n1 20.689
R21329 a_3152_n45.n0 a_3152_n45.t2 362.857
R21330 a_3152_n45.t4 a_3152_n45.t3 337.399
R21331 a_3152_n45.t3 a_3152_n45.t5 298.839
R21332 a_3152_n45.n0 a_3152_n45.t4 280.405
R21333 a_3152_n45.n1 a_3152_n45.t0 200
R21334 a_3152_n45.n1 a_3152_n45.n0 172.311
R21335 a_3152_n45.n2 a_3152_n45.n1 24
R21336 a_3152_n45.n1 a_3152_n45.t1 21.212
R21337 a_852_n286.n0 a_852_n286.t1 362.857
R21338 a_852_n286.t3 a_852_n286.t4 337.399
R21339 a_852_n286.t4 a_852_n286.t5 298.839
R21340 a_852_n286.n0 a_852_n286.t3 280.405
R21341 a_852_n286.n1 a_852_n286.t0 200
R21342 a_852_n286.n1 a_852_n286.n0 172.311
R21343 a_852_n286.n2 a_852_n286.n1 24
R21344 a_852_n286.n1 a_852_n286.t2 21.212
R21345 a_947_n271.n0 a_947_n271.t1 358.166
R21346 a_947_n271.t4 a_947_n271.t5 337.399
R21347 a_947_n271.t5 a_947_n271.t3 285.986
R21348 a_947_n271.n0 a_947_n271.t4 282.573
R21349 a_947_n271.n1 a_947_n271.t2 202.857
R21350 a_947_n271.n1 a_947_n271.n0 173.817
R21351 a_947_n271.n1 a_947_n271.t0 20.826
R21352 a_947_n271.n2 a_947_n271.n1 20.689
R21353 a_8327_437.n0 a_8327_437.t2 362.857
R21354 a_8327_437.t4 a_8327_437.t3 337.399
R21355 a_8327_437.t3 a_8327_437.t5 298.839
R21356 a_8327_437.n0 a_8327_437.t4 280.405
R21357 a_8327_437.n1 a_8327_437.t0 200
R21358 a_8327_437.n1 a_8327_437.n0 172.311
R21359 a_8327_437.n2 a_8327_437.n1 24
R21360 a_8327_437.n1 a_8327_437.t1 21.212
R21361 a_8422_452.n0 a_8422_452.t1 358.166
R21362 a_8422_452.t5 a_8422_452.t4 337.399
R21363 a_8422_452.t4 a_8422_452.t3 285.986
R21364 a_8422_452.n0 a_8422_452.t5 282.573
R21365 a_8422_452.n1 a_8422_452.t2 202.857
R21366 a_8422_452.n1 a_8422_452.n0 173.817
R21367 a_8422_452.n1 a_8422_452.t0 20.826
R21368 a_8422_452.n2 a_8422_452.n1 20.689
R21369 a_1522_1698.n0 a_1522_1698.t1 358.166
R21370 a_1522_1698.t3 a_1522_1698.t5 337.399
R21371 a_1522_1698.t5 a_1522_1698.t4 285.986
R21372 a_1522_1698.n0 a_1522_1698.t3 282.573
R21373 a_1522_1698.n1 a_1522_1698.t2 202.857
R21374 a_1522_1698.n1 a_1522_1698.n0 173.817
R21375 a_1522_1698.n1 a_1522_1698.t0 20.826
R21376 a_1522_1698.n2 a_1522_1698.n1 20.689
R21377 a_6040_693.t0 a_6040_693.t1 242.857
R21378 a_8915_n1053.t0 a_8915_n1053.t1 242.857
R21379 a_865_3666.t0 a_865_3666.t1 242.857
R21380 a_3165_2180.t0 a_3165_2180.t1 242.857
R21381 SA_OUT[11].n1 SA_OUT[11].t3 661.027
R21382 SA_OUT[11].n1 SA_OUT[11].t4 392.255
R21383 SA_OUT[11].n2 SA_OUT[11].t1 223.716
R21384 SA_OUT[11].n0 SA_OUT[11].t2 153.977
R21385 SA_OUT[11].n2 SA_OUT[11].n1 143.764
R21386 SA_OUT[11].n0 SA_OUT[11].t0 59.86
R21387 SA_OUT[11] SA_OUT[11].n3 14.218
R21388 SA_OUT[11].n3 SA_OUT[11].n0 3.764
R21389 SA_OUT[11].n3 SA_OUT[11].n2 0.752
R21390 a_6635_n1371.n1 a_6635_n1371.t4 550.94
R21391 a_6635_n1371.n1 a_6635_n1371.t3 500.621
R21392 a_6635_n1371.t2 a_6635_n1371.n2 192.787
R21393 a_6635_n1371.n0 a_6635_n1371.t0 163.997
R21394 a_6635_n1371.n2 a_6635_n1371.n1 149.035
R21395 a_6635_n1371.n0 a_6635_n1371.t1 54.068
R21396 a_6635_n1371.n2 a_6635_n1371.n0 17.317
R21397 a_6727_n1770.t0 a_6727_n1770.n0 182.779
R21398 a_6727_n1770.n0 a_6727_n1770.t1 111.474
R21399 a_2015_4148.t0 a_2015_4148.t1 242.857
R21400 a_4972_693.n0 a_4972_693.t2 358.166
R21401 a_4972_693.t4 a_4972_693.t3 337.399
R21402 a_4972_693.t3 a_4972_693.t5 285.986
R21403 a_4972_693.n0 a_4972_693.t4 282.573
R21404 a_4972_693.n1 a_4972_693.t0 202.857
R21405 a_4972_693.n1 a_4972_693.n0 173.817
R21406 a_4972_693.n1 a_4972_693.t1 20.826
R21407 a_4972_693.n2 a_4972_693.n1 20.689
R21408 a_4877_678.n0 a_4877_678.t1 362.857
R21409 a_4877_678.t5 a_4877_678.t4 337.399
R21410 a_4877_678.t4 a_4877_678.t3 298.839
R21411 a_4877_678.n0 a_4877_678.t5 280.405
R21412 a_4877_678.n1 a_4877_678.t2 200
R21413 a_4877_678.n1 a_4877_678.n0 172.311
R21414 a_4877_678.n2 a_4877_678.n1 24
R21415 a_4877_678.n1 a_4877_678.t0 21.212
R21416 a_4397_3666.n0 a_4397_3666.t1 358.166
R21417 a_4397_3666.t4 a_4397_3666.t5 337.399
R21418 a_4397_3666.t5 a_4397_3666.t3 285.986
R21419 a_4397_3666.n0 a_4397_3666.t4 282.573
R21420 a_4397_3666.n1 a_4397_3666.t2 202.857
R21421 a_4397_3666.n1 a_4397_3666.n0 173.817
R21422 a_4397_3666.n1 a_4397_3666.t0 20.826
R21423 a_4397_3666.n2 a_4397_3666.n1 20.689
R21424 a_4767_3666.t0 a_4767_3666.t1 242.857
R21425 a_5452_1924.n0 a_5452_1924.t1 362.857
R21426 a_5452_1924.t3 a_5452_1924.t4 337.399
R21427 a_5452_1924.t4 a_5452_1924.t5 298.839
R21428 a_5452_1924.n0 a_5452_1924.t3 280.405
R21429 a_5452_1924.n1 a_5452_1924.t0 200
R21430 a_5452_1924.n1 a_5452_1924.n0 172.311
R21431 a_5452_1924.n2 a_5452_1924.n1 24
R21432 a_5452_1924.n1 a_5452_1924.t2 21.212
R21433 a_2652_n2234.n2 a_2652_n2234.t0 282.97
R21434 a_2652_n2234.n1 a_2652_n2234.t4 240.683
R21435 a_2652_n2234.n0 a_2652_n2234.t2 209.208
R21436 a_2652_n2234.n0 a_2652_n2234.t3 194.167
R21437 a_2652_n2234.t1 a_2652_n2234.n2 183.404
R21438 a_2652_n2234.n1 a_2652_n2234.n0 14.805
R21439 a_2652_n2234.n2 a_2652_n2234.n1 6.415
R21440 a_2775_n2132.n0 a_2775_n2132.t2 489.336
R21441 a_2775_n2132.n0 a_2775_n2132.t1 243.258
R21442 a_2775_n2132.t0 a_2775_n2132.n0 214.415
R21443 a_1522_n812.n0 a_1522_n812.t2 358.166
R21444 a_1522_n812.t3 a_1522_n812.t5 337.399
R21445 a_1522_n812.t5 a_1522_n812.t4 285.986
R21446 a_1522_n812.n0 a_1522_n812.t3 282.573
R21447 a_1522_n812.n1 a_1522_n812.t0 202.857
R21448 a_1522_n812.n1 a_1522_n812.n0 173.817
R21449 a_1522_n812.n1 a_1522_n812.t1 20.826
R21450 a_1522_n812.n2 a_1522_n812.n1 20.689
R21451 a_742_1939.t0 a_742_1939.t1 242.857
R21452 a_8792_452.t0 a_8792_452.t1 242.857
R21453 a_4397_n512.n0 a_4397_n512.t1 358.166
R21454 a_4397_n512.t5 a_4397_n512.t3 337.399
R21455 a_4397_n512.t3 a_4397_n512.t4 285.986
R21456 a_4397_n512.n0 a_4397_n512.t5 282.573
R21457 a_4397_n512.n1 a_4397_n512.t0 202.857
R21458 a_4397_n512.n1 a_4397_n512.n0 173.817
R21459 a_4397_n512.n1 a_4397_n512.t2 20.826
R21460 a_4397_n512.n2 a_4397_n512.n1 20.689
R21461 a_4302_n527.n0 a_4302_n527.t1 362.857
R21462 a_4302_n527.t3 a_4302_n527.t5 337.399
R21463 a_4302_n527.t5 a_4302_n527.t4 298.839
R21464 a_4302_n527.n0 a_4302_n527.t3 280.405
R21465 a_4302_n527.n1 a_4302_n527.t2 200
R21466 a_4302_n527.n1 a_4302_n527.n0 172.311
R21467 a_4302_n527.n2 a_4302_n527.n1 24
R21468 a_4302_n527.n1 a_4302_n527.t0 21.212
R21469 a_4890_4686.t0 a_4890_4686.t1 242.857
R21470 a_1317_3184.t0 a_1317_3184.t1 242.857
R21471 a_5547_1216.n0 a_5547_1216.t1 358.166
R21472 a_5547_1216.t5 a_5547_1216.t3 337.399
R21473 a_5547_1216.t3 a_5547_1216.t4 285.986
R21474 a_5547_1216.n0 a_5547_1216.t5 282.573
R21475 a_5547_1216.n1 a_5547_1216.t0 202.857
R21476 a_5547_1216.n1 a_5547_1216.n0 173.817
R21477 a_5547_1216.n1 a_5547_1216.t2 20.826
R21478 a_5547_1216.n2 a_5547_1216.n1 20.689
R21479 a_5452_1201.n0 a_5452_1201.t2 362.857
R21480 a_5452_1201.t3 a_5452_1201.t4 337.399
R21481 a_5452_1201.t4 a_5452_1201.t5 298.839
R21482 a_5452_1201.n0 a_5452_1201.t3 280.405
R21483 a_5452_1201.n1 a_5452_1201.t0 200
R21484 a_5452_1201.n1 a_5452_1201.n0 172.311
R21485 a_5452_1201.n2 a_5452_1201.n1 24
R21486 a_5452_1201.n1 a_5452_1201.t1 21.212
R21487 a_290_4445.t0 a_290_4445.t1 242.857
R21488 a_n2677_n5092.t0 a_n2677_n5092.t1 42.705
R21489 a_4192_4445.t0 a_4192_4445.t1 242.857
R21490 a_6122_n812.n0 a_6122_n812.t2 358.166
R21491 a_6122_n812.t4 a_6122_n812.t3 337.399
R21492 a_6122_n812.t3 a_6122_n812.t5 285.986
R21493 a_6122_n812.n0 a_6122_n812.t4 282.573
R21494 a_6122_n812.n1 a_6122_n812.t0 202.857
R21495 a_6122_n812.n1 a_6122_n812.n0 173.817
R21496 a_6122_n812.n1 a_6122_n812.t1 20.826
R21497 a_6122_n812.n2 a_6122_n812.n1 20.689
R21498 a_3740_n812.t0 a_3740_n812.t1 242.857
R21499 a_3042_1457.t0 a_3042_1457.t1 242.857
R21500 a_13602_n5092.t0 a_13602_n5092.t1 42.705
R21501 a_13637_n5293.n0 a_13637_n5293.t0 65.063
R21502 a_13637_n5293.n0 a_13637_n5293.t2 42.011
R21503 a_13637_n5293.t1 a_13637_n5293.n0 2.113
R21504 a_5465_4445.t0 a_5465_4445.t1 242.857
R21505 a_8327_4430.n0 a_8327_4430.t1 362.857
R21506 a_8327_4430.t5 a_8327_4430.t3 337.399
R21507 a_8327_4430.t3 a_8327_4430.t4 298.839
R21508 a_8327_4430.n0 a_8327_4430.t5 280.405
R21509 a_8327_4430.n1 a_8327_4430.t2 200
R21510 a_8327_4430.n1 a_8327_4430.n0 172.311
R21511 a_8327_4430.n2 a_8327_4430.n1 24
R21512 a_8327_4430.n1 a_8327_4430.t0 21.212
R21513 a_4397_n271.n0 a_4397_n271.t1 358.166
R21514 a_4397_n271.t4 a_4397_n271.t5 337.399
R21515 a_4397_n271.t5 a_4397_n271.t3 285.986
R21516 a_4397_n271.n0 a_4397_n271.t4 282.573
R21517 a_4397_n271.n1 a_4397_n271.t2 202.857
R21518 a_4397_n271.n1 a_4397_n271.n0 173.817
R21519 a_4397_n271.n1 a_4397_n271.t0 20.826
R21520 a_4397_n271.n2 a_4397_n271.n1 20.689
R21521 a_8217_4686.t0 a_8217_4686.t1 242.857
R21522 a_6615_2180.t0 a_6615_2180.t1 242.857
R21523 a_867_n4378.n3 a_867_n4378.t3 475.39
R21524 a_867_n4378.n3 a_867_n4378.n2 306.026
R21525 a_867_n4378.t4 a_867_n4378.t6 228.696
R21526 a_867_n4378.n2 a_867_n4378.t1 185.704
R21527 a_867_n4378.n0 a_867_n4378.t4 126.761
R21528 a_867_n4378.n1 a_867_n4378.t5 126.284
R21529 a_867_n4378.n1 a_867_n4378.t0 126.284
R21530 a_867_n4378.t2 a_867_n4378.n3 124.375
R21531 a_867_n4378.t0 a_867_n4378.n0 115.122
R21532 a_867_n4378.n0 a_867_n4378.t7 111.229
R21533 a_867_n4378.n2 a_867_n4378.n1 8.764
R21534 a_867_n6849.t0 a_867_n6849.t1 42.707
R21535 a_1522_1216.n0 a_1522_1216.t2 358.166
R21536 a_1522_1216.t3 a_1522_1216.t5 337.399
R21537 a_1522_1216.t5 a_1522_1216.t4 285.986
R21538 a_1522_1216.n0 a_1522_1216.t3 282.573
R21539 a_1522_1216.n1 a_1522_1216.t0 202.857
R21540 a_1522_1216.n1 a_1522_1216.n0 173.817
R21541 a_1522_1216.n1 a_1522_1216.t1 20.826
R21542 a_1522_1216.n2 a_1522_1216.n1 20.689
R21543 a_6027_n45.n0 a_6027_n45.t2 362.857
R21544 a_6027_n45.t4 a_6027_n45.t3 337.399
R21545 a_6027_n45.t3 a_6027_n45.t5 298.839
R21546 a_6027_n45.n0 a_6027_n45.t4 280.405
R21547 a_6027_n45.n1 a_6027_n45.t0 200
R21548 a_6027_n45.n1 a_6027_n45.n0 172.311
R21549 a_6027_n45.n2 a_6027_n45.n1 24
R21550 a_6027_n45.n1 a_6027_n45.t1 21.212
R21551 a_2590_452.t0 a_2590_452.t1 242.857
R21552 a_6027_1442.n0 a_6027_1442.t0 362.857
R21553 a_6027_1442.t3 a_6027_1442.t4 337.399
R21554 a_6027_1442.t4 a_6027_1442.t5 298.839
R21555 a_6027_1442.n0 a_6027_1442.t3 280.405
R21556 a_6027_1442.n1 a_6027_1442.t2 200
R21557 a_6027_1442.n1 a_6027_1442.n0 172.311
R21558 a_6027_1442.n2 a_6027_1442.n1 24
R21559 a_6027_1442.n1 a_6027_1442.t1 21.212
R21560 a_5342_693.t0 a_5342_693.t1 242.857
R21561 a_6812_n5293.n0 a_6812_n5293.t0 65.063
R21562 a_6812_n5293.n0 a_6812_n5293.t2 42.011
R21563 a_6812_n5293.t1 a_6812_n5293.n0 2.113
R21564 a_2590_n512.t0 a_2590_n512.t1 242.857
R21565 a_4972_3907.n0 a_4972_3907.t1 358.166
R21566 a_4972_3907.t3 a_4972_3907.t5 337.399
R21567 a_4972_3907.t5 a_4972_3907.t4 285.986
R21568 a_4972_3907.n0 a_4972_3907.t3 282.573
R21569 a_4972_3907.n1 a_4972_3907.t2 202.857
R21570 a_4972_3907.n1 a_4972_3907.n0 173.817
R21571 a_4972_3907.n1 a_4972_3907.t0 20.826
R21572 a_4972_3907.n2 a_4972_3907.n1 20.689
R21573 a_4877_3892.n0 a_4877_3892.t1 362.857
R21574 a_4877_3892.t4 a_4877_3892.t3 337.399
R21575 a_4877_3892.t3 a_4877_3892.t5 298.839
R21576 a_4877_3892.n0 a_4877_3892.t4 280.405
R21577 a_4877_3892.n1 a_4877_3892.t2 200
R21578 a_4877_3892.n1 a_4877_3892.n0 172.311
R21579 a_4877_3892.n2 a_4877_3892.n1 24
R21580 a_4877_3892.n1 a_4877_3892.t0 21.212
R21581 a_277_2928.n0 a_277_2928.t2 362.857
R21582 a_277_2928.t3 a_277_2928.t4 337.399
R21583 a_277_2928.t4 a_277_2928.t5 298.839
R21584 a_277_2928.n0 a_277_2928.t3 280.405
R21585 a_277_2928.n1 a_277_2928.t0 200
R21586 a_277_2928.n1 a_277_2928.n0 172.311
R21587 a_277_2928.n2 a_277_2928.n1 24
R21588 a_277_2928.n1 a_277_2928.t1 21.212
R21589 a_7642_4445.t0 a_7642_4445.t1 242.857
R21590 a_8997_3907.n0 a_8997_3907.t1 358.166
R21591 a_8997_3907.t4 a_8997_3907.t5 337.399
R21592 a_8997_3907.t5 a_8997_3907.t3 285.986
R21593 a_8997_3907.n0 a_8997_3907.t4 282.573
R21594 a_8997_3907.n1 a_8997_3907.t2 202.857
R21595 a_8997_3907.n1 a_8997_3907.n0 173.817
R21596 a_8997_3907.n1 a_8997_3907.t0 20.826
R21597 a_8997_3907.n2 a_8997_3907.n1 20.689
R21598 a_9367_3907.t0 a_9367_3907.t1 242.857
R21599 a_3822_2662.n0 a_3822_2662.t1 358.166
R21600 a_3822_2662.t5 a_3822_2662.t4 337.399
R21601 a_3822_2662.t4 a_3822_2662.t3 285.986
R21602 a_3822_2662.n0 a_3822_2662.t5 282.573
R21603 a_3822_2662.n1 a_3822_2662.t2 202.857
R21604 a_3822_2662.n1 a_3822_2662.n0 173.817
R21605 a_3822_2662.n1 a_3822_2662.t0 20.826
R21606 a_3822_2662.n2 a_3822_2662.n1 20.689
R21607 a_1168_n2086.t0 a_1168_n2086.t1 34.8
R21608 a_6122_n1053.n0 a_6122_n1053.t1 358.166
R21609 a_6122_n1053.t3 a_6122_n1053.t5 337.399
R21610 a_6122_n1053.t5 a_6122_n1053.t4 285.986
R21611 a_6122_n1053.n0 a_6122_n1053.t3 282.573
R21612 a_6122_n1053.n1 a_6122_n1053.t0 202.857
R21613 a_6122_n1053.n1 a_6122_n1053.n0 173.817
R21614 a_6122_n1053.n1 a_6122_n1053.t2 20.826
R21615 a_6122_n1053.n2 a_6122_n1053.n1 20.689
R21616 a_6027_n1068.n0 a_6027_n1068.t1 362.857
R21617 a_6027_n1068.t3 a_6027_n1068.t4 337.399
R21618 a_6027_n1068.t4 a_6027_n1068.t5 298.839
R21619 a_6027_n1068.n0 a_6027_n1068.t3 280.405
R21620 a_6027_n1068.n1 a_6027_n1068.t2 200
R21621 a_6027_n1068.n1 a_6027_n1068.n0 172.311
R21622 a_6027_n1068.n2 a_6027_n1068.n1 24
R21623 a_6027_n1068.n1 a_6027_n1068.t0 21.212
R21624 a_1427_4430.n0 a_1427_4430.t0 362.857
R21625 a_1427_4430.t3 a_1427_4430.t4 337.399
R21626 a_1427_4430.t4 a_1427_4430.t5 298.839
R21627 a_1427_4430.n0 a_1427_4430.t3 280.405
R21628 a_1427_4430.n1 a_1427_4430.t2 200
R21629 a_1427_4430.n1 a_1427_4430.n0 172.311
R21630 a_1427_4430.n2 a_1427_4430.n1 24
R21631 a_1427_4430.n1 a_1427_4430.t1 21.212
R21632 a_3165_3184.t0 a_3165_3184.t1 242.857
R21633 a_6027_3169.n0 a_6027_3169.t2 362.857
R21634 a_6027_3169.t5 a_6027_3169.t3 337.399
R21635 a_6027_3169.t3 a_6027_3169.t4 298.839
R21636 a_6027_3169.n0 a_6027_3169.t5 280.405
R21637 a_6027_3169.n1 a_6027_3169.t0 200
R21638 a_6027_3169.n1 a_6027_3169.n0 172.311
R21639 a_6027_3169.n2 a_6027_3169.n1 24
R21640 a_6027_3169.n1 a_6027_3169.t1 21.212
R21641 a_7067_975.t0 a_7067_975.t1 242.857
R21642 a_8915_4445.t0 a_8915_4445.t1 242.857
R21643 a_7765_975.t0 a_7765_975.t1 242.857
R21644 a_2097_452.n0 a_2097_452.t0 358.166
R21645 a_2097_452.t5 a_2097_452.t4 337.399
R21646 a_2097_452.t4 a_2097_452.t3 285.986
R21647 a_2097_452.n0 a_2097_452.t5 282.573
R21648 a_2097_452.n1 a_2097_452.t2 202.857
R21649 a_2097_452.n1 a_2097_452.n0 173.817
R21650 a_2097_452.n1 a_2097_452.t1 20.826
R21651 a_2097_452.n2 a_2097_452.n1 20.689
R21652 a_2467_452.t0 a_2467_452.t1 242.857
R21653 a_3727_437.n0 a_3727_437.t1 362.857
R21654 a_3727_437.t4 a_3727_437.t3 337.399
R21655 a_3727_437.t3 a_3727_437.t5 298.839
R21656 a_3727_437.n0 a_3727_437.t4 280.405
R21657 a_3727_437.n1 a_3727_437.t2 200
R21658 a_3727_437.n1 a_3727_437.n0 172.311
R21659 a_3727_437.n2 a_3727_437.n1 24
R21660 a_3727_437.n1 a_3727_437.t0 21.212
R21661 a_3822_452.n0 a_3822_452.t2 358.166
R21662 a_3822_452.t4 a_3822_452.t3 337.399
R21663 a_3822_452.t3 a_3822_452.t5 285.986
R21664 a_3822_452.n0 a_3822_452.t4 282.573
R21665 a_3822_452.n1 a_3822_452.t0 202.857
R21666 a_3822_452.n1 a_3822_452.n0 173.817
R21667 a_3822_452.n1 a_3822_452.t1 20.826
R21668 a_3822_452.n2 a_3822_452.n1 20.689
R21669 a_5452_n1068.n0 a_5452_n1068.t1 362.857
R21670 a_5452_n1068.t5 a_5452_n1068.t3 337.399
R21671 a_5452_n1068.t3 a_5452_n1068.t4 298.839
R21672 a_5452_n1068.n0 a_5452_n1068.t5 280.405
R21673 a_5452_n1068.n1 a_5452_n1068.t0 200
R21674 a_5452_n1068.n1 a_5452_n1068.n0 172.311
R21675 a_5452_n1068.n2 a_5452_n1068.n1 24
R21676 a_5452_n1068.n1 a_5452_n1068.t2 21.212
R21677 a_852_960.n0 a_852_960.t2 362.857
R21678 a_852_960.t3 a_852_960.t5 337.399
R21679 a_852_960.t5 a_852_960.t4 298.839
R21680 a_852_960.n0 a_852_960.t3 280.405
R21681 a_852_960.n1 a_852_960.t0 200
R21682 a_852_960.n1 a_852_960.n0 172.311
R21683 a_852_960.n2 a_852_960.n1 24
R21684 a_852_960.n1 a_852_960.t1 21.212
R21685 a_1440_693.t0 a_1440_693.t1 242.857
R21686 a_6040_4148.t0 a_6040_4148.t1 242.857
R21687 a_7190_2180.t0 a_7190_2180.t1 242.857
R21688 a_5547_4445.n0 a_5547_4445.t0 358.166
R21689 a_5547_4445.t5 a_5547_4445.t3 337.399
R21690 a_5547_4445.t3 a_5547_4445.t4 285.986
R21691 a_5547_4445.n0 a_5547_4445.t5 282.573
R21692 a_5547_4445.n1 a_5547_4445.t2 202.857
R21693 a_5547_4445.n1 a_5547_4445.n0 173.817
R21694 a_5547_4445.n1 a_5547_4445.t1 20.826
R21695 a_5547_4445.n2 a_5547_4445.n1 20.689
R21696 a_5452_4430.n0 a_5452_4430.t2 362.857
R21697 a_5452_4430.t3 a_5452_4430.t4 337.399
R21698 a_5452_4430.t4 a_5452_4430.t5 298.839
R21699 a_5452_4430.n0 a_5452_4430.t3 280.405
R21700 a_5452_4430.n1 a_5452_4430.t0 200
R21701 a_5452_4430.n1 a_5452_4430.n0 172.311
R21702 a_5452_4430.n2 a_5452_4430.n1 24
R21703 a_5452_4430.n1 a_5452_4430.t1 21.212
R21704 a_8792_3666.t0 a_8792_3666.t1 242.857
R21705 a_4043_n2086.t0 a_4043_n2086.t1 34.8
R21706 a_2590_2943.t0 a_2590_2943.t1 242.857
R21707 a_4972_n271.n0 a_4972_n271.t1 358.166
R21708 a_4972_n271.t3 a_4972_n271.t5 337.399
R21709 a_4972_n271.t5 a_4972_n271.t4 285.986
R21710 a_4972_n271.n0 a_4972_n271.t3 282.573
R21711 a_4972_n271.n1 a_4972_n271.t2 202.857
R21712 a_4972_n271.n1 a_4972_n271.n0 173.817
R21713 a_4972_n271.n1 a_4972_n271.t0 20.826
R21714 a_4972_n271.n2 a_4972_n271.n1 20.689
R21715 a_8422_n512.n0 a_8422_n512.t2 358.166
R21716 a_8422_n512.t4 a_8422_n512.t3 337.399
R21717 a_8422_n512.t3 a_8422_n512.t5 285.986
R21718 a_8422_n512.n0 a_8422_n512.t4 282.573
R21719 a_8422_n512.n1 a_8422_n512.t0 202.857
R21720 a_8422_n512.n1 a_8422_n512.n0 173.817
R21721 a_8422_n512.n1 a_8422_n512.t1 20.826
R21722 a_8422_n512.n2 a_8422_n512.n1 20.689
R21723 a_2467_4148.t0 a_2467_4148.t1 242.857
R21724 a_5342_3184.t0 a_5342_3184.t1 242.857
R21725 a_8997_n271.n0 a_8997_n271.t2 358.166
R21726 a_8997_n271.t4 a_8997_n271.t5 337.399
R21727 a_8997_n271.t5 a_8997_n271.t3 285.986
R21728 a_8997_n271.n0 a_8997_n271.t4 282.573
R21729 a_8997_n271.n1 a_8997_n271.t0 202.857
R21730 a_8997_n271.n1 a_8997_n271.n0 173.817
R21731 a_8997_n271.n1 a_8997_n271.t1 20.826
R21732 a_8997_n271.n2 a_8997_n271.n1 20.689
R21733 a_9367_n271.t0 a_9367_n271.t1 242.857
R21734 a_2085_n1770.n0 a_2085_n1770.t1 325.682
R21735 a_2085_n1770.n0 a_2085_n1770.t2 322.294
R21736 a_2085_n1770.t0 a_2085_n1770.n0 73.623
R21737 a_360_n1770.n0 a_360_n1770.t2 322.294
R21738 a_360_n1770.n1 a_360_n1770.n0 229.466
R21739 a_360_n1770.t0 a_360_n1770.n1 151.15
R21740 a_360_n1770.n0 a_360_n1770.t1 73.623
R21741 a_402_n1770.t0 a_402_n1770.n0 182.779
R21742 a_402_n1770.n0 a_402_n1770.t1 111.474
R21743 a_3042_4686.t0 a_3042_4686.t1 242.857
R21744 a_4972_3425.n0 a_4972_3425.t2 358.166
R21745 a_4972_3425.t3 a_4972_3425.t5 337.399
R21746 a_4972_3425.t5 a_4972_3425.t4 285.986
R21747 a_4972_3425.n0 a_4972_3425.t3 282.573
R21748 a_4972_3425.n1 a_4972_3425.t0 202.857
R21749 a_4972_3425.n1 a_4972_3425.n0 173.817
R21750 a_4972_3425.n1 a_4972_3425.t1 20.826
R21751 a_4972_3425.n2 a_4972_3425.n1 20.689
R21752 a_4877_3410.n0 a_4877_3410.t2 362.857
R21753 a_4877_3410.t4 a_4877_3410.t3 337.399
R21754 a_4877_3410.t3 a_4877_3410.t5 298.839
R21755 a_4877_3410.n0 a_4877_3410.t4 280.405
R21756 a_4877_3410.n1 a_4877_3410.t0 200
R21757 a_4877_3410.n1 a_4877_3410.n0 172.311
R21758 a_4877_3410.n2 a_4877_3410.n1 24
R21759 a_4877_3410.n1 a_4877_3410.t1 21.212
R21760 a_6122_1457.n0 a_6122_1457.t1 358.166
R21761 a_6122_1457.t3 a_6122_1457.t5 337.399
R21762 a_6122_1457.t5 a_6122_1457.t4 285.986
R21763 a_6122_1457.n0 a_6122_1457.t3 282.573
R21764 a_6122_1457.n1 a_6122_1457.t2 202.857
R21765 a_6122_1457.n1 a_6122_1457.n0 173.817
R21766 a_6122_1457.n1 a_6122_1457.t0 20.826
R21767 a_6122_1457.n2 a_6122_1457.n1 20.689
R21768 a_1440_2180.t0 a_1440_2180.t1 242.857
R21769 a_6615_3184.t0 a_6615_3184.t1 242.857
R21770 a_8327_n1068.n0 a_8327_n1068.t1 362.857
R21771 a_8327_n1068.t5 a_8327_n1068.t3 337.399
R21772 a_8327_n1068.t3 a_8327_n1068.t4 298.839
R21773 a_8327_n1068.n0 a_8327_n1068.t5 280.405
R21774 a_8327_n1068.n1 a_8327_n1068.t0 200
R21775 a_8327_n1068.n1 a_8327_n1068.n0 172.311
R21776 a_8327_n1068.n2 a_8327_n1068.n1 24
R21777 a_8327_n1068.n1 a_8327_n1068.t2 21.212
R21778 a_8997_3425.n0 a_8997_3425.t2 358.166
R21779 a_8997_3425.t4 a_8997_3425.t5 337.399
R21780 a_8997_3425.t5 a_8997_3425.t3 285.986
R21781 a_8997_3425.n0 a_8997_3425.t4 282.573
R21782 a_8997_3425.n1 a_8997_3425.t0 202.857
R21783 a_8997_3425.n1 a_8997_3425.n0 173.817
R21784 a_8997_3425.n1 a_8997_3425.t1 20.826
R21785 a_8997_3425.n2 a_8997_3425.n1 20.689
R21786 a_9367_3425.t0 a_9367_3425.t1 242.857
R21787 a_6602_678.n0 a_6602_678.t1 362.857
R21788 a_6602_678.t3 a_6602_678.t5 337.399
R21789 a_6602_678.t5 a_6602_678.t4 298.839
R21790 a_6602_678.n0 a_6602_678.t3 280.405
R21791 a_6602_678.n1 a_6602_678.t2 200
R21792 a_6602_678.n1 a_6602_678.n0 172.311
R21793 a_6602_678.n2 a_6602_678.n1 24
R21794 a_6602_678.n1 a_6602_678.t0 21.212
R21795 a_6697_693.n0 a_6697_693.t2 358.166
R21796 a_6697_693.t4 a_6697_693.t3 337.399
R21797 a_6697_693.t3 a_6697_693.t5 285.986
R21798 a_6697_693.n0 a_6697_693.t4 282.573
R21799 a_6697_693.n1 a_6697_693.t0 202.857
R21800 a_6697_693.n1 a_6697_693.n0 173.817
R21801 a_6697_693.n1 a_6697_693.t1 20.826
R21802 a_6697_693.n2 a_6697_693.n1 20.689
R21803 a_4745_n7203.n0 a_4745_n7203.t0 63.08
R21804 a_4745_n7203.t1 a_4745_n7203.n0 41.306
R21805 a_4745_n7203.n0 a_4745_n7203.t2 2.251
R21806 a_18_n7203.n0 a_18_n7203.t0 63.08
R21807 a_18_n7203.n0 a_18_n7203.t2 41.305
R21808 a_18_n7203.t1 a_18_n7203.n0 2.251
R21809 a_3617_2421.t0 a_3617_2421.t1 242.857
R21810 a_2318_n2086.t0 a_2318_n2086.t1 34.8
R21811 a_1522_4445.n0 a_1522_4445.t2 358.166
R21812 a_1522_4445.t3 a_1522_4445.t5 337.399
R21813 a_1522_4445.t5 a_1522_4445.t4 285.986
R21814 a_1522_4445.n0 a_1522_4445.t3 282.573
R21815 a_1522_4445.n1 a_1522_4445.t0 202.857
R21816 a_1522_4445.n1 a_1522_4445.n0 173.817
R21817 a_1522_4445.n1 a_1522_4445.t1 20.826
R21818 a_1522_4445.n2 a_1522_4445.n1 20.689
R21819 a_3617_n271.t0 a_3617_n271.t1 242.857
R21820 a_6027_4671.n0 a_6027_4671.t2 362.857
R21821 a_6027_4671.t3 a_6027_4671.t4 337.399
R21822 a_6027_4671.t4 a_6027_4671.t5 298.839
R21823 a_6027_4671.n0 a_6027_4671.t3 280.405
R21824 a_6027_4671.n1 a_6027_4671.t0 200
R21825 a_6027_4671.n1 a_6027_4671.n0 172.311
R21826 a_6027_4671.n2 a_6027_4671.n1 24
R21827 a_6027_4671.n1 a_6027_4671.t1 21.212
R21828 a_3247_3184.n0 a_3247_3184.t0 358.166
R21829 a_3247_3184.t5 a_3247_3184.t3 337.399
R21830 a_3247_3184.t3 a_3247_3184.t4 285.986
R21831 a_3247_3184.n0 a_3247_3184.t5 282.573
R21832 a_3247_3184.n1 a_3247_3184.t1 202.857
R21833 a_3247_3184.n1 a_3247_3184.n0 173.817
R21834 a_3247_3184.n1 a_3247_3184.t2 20.826
R21835 a_3247_3184.n2 a_3247_3184.n1 20.689
R21836 a_3152_3169.n0 a_3152_3169.t2 362.857
R21837 a_3152_3169.t3 a_3152_3169.t4 337.399
R21838 a_3152_3169.t4 a_3152_3169.t5 298.839
R21839 a_3152_3169.n0 a_3152_3169.t3 280.405
R21840 a_3152_3169.n1 a_3152_3169.t0 200
R21841 a_3152_3169.n1 a_3152_3169.n0 172.311
R21842 a_3152_3169.n2 a_3152_3169.n1 24
R21843 a_3152_3169.n1 a_3152_3169.t1 21.212
R21844 a_2015_1939.t0 a_2015_1939.t1 242.857
R21845 ADC14_OUT[2].n0 ADC14_OUT[2].t4 1354.27
R21846 ADC14_OUT[2].n0 ADC14_OUT[2].t3 821.954
R21847 ADC14_OUT[2].n3 ADC14_OUT[2].t0 338.856
R21848 ADC14_OUT[2].n2 ADC14_OUT[2].t1 266.575
R21849 ADC14_OUT[2].n1 ADC14_OUT[2].n0 149.035
R21850 ADC14_OUT[2].n1 ADC14_OUT[2].t2 46.723
R21851 ADC14_OUT[2].n3 ADC14_OUT[2].n2 45.176
R21852 ADC14_OUT[2] ADC14_OUT[2].n3 37.985
R21853 ADC14_OUT[2].n2 ADC14_OUT[2].n1 17.317
R21854 a_1427_n45.n0 a_1427_n45.t0 362.857
R21855 a_1427_n45.t4 a_1427_n45.t3 337.399
R21856 a_1427_n45.t3 a_1427_n45.t5 298.839
R21857 a_1427_n45.n0 a_1427_n45.t4 280.405
R21858 a_1427_n45.n1 a_1427_n45.t2 200
R21859 a_1427_n45.n1 a_1427_n45.n0 172.311
R21860 a_1427_n45.n2 a_1427_n45.n1 24
R21861 a_1427_n45.n1 a_1427_n45.t1 21.212
R21862 ADC4_OUT[1].n0 ADC4_OUT[1].t4 1355.37
R21863 ADC4_OUT[1].n0 ADC4_OUT[1].t3 820.859
R21864 ADC4_OUT[1].n3 ADC4_OUT[1].t0 326.879
R21865 ADC4_OUT[1].n2 ADC4_OUT[1].t1 266.644
R21866 ADC4_OUT[1].n1 ADC4_OUT[1].n0 149.035
R21867 ADC4_OUT[1].n3 ADC4_OUT[1].n2 57.223
R21868 ADC4_OUT[1].n1 ADC4_OUT[1].t2 45.968
R21869 ADC4_OUT[1] ADC4_OUT[1].n3 45.847
R21870 ADC4_OUT[1].n2 ADC4_OUT[1].n1 17.317
R21871 a_1129_n5850.n0 a_1129_n5850.t4 1465.51
R21872 a_1129_n5850.n0 a_1129_n5850.t3 712.44
R21873 a_1129_n5850.n1 a_1129_n5850.t0 375.067
R21874 a_1129_n5850.n1 a_1129_n5850.t1 272.668
R21875 a_1129_n5850.n2 a_1129_n5850.n0 143.764
R21876 a_1129_n5850.t2 a_1129_n5850.n2 78.193
R21877 a_1129_n5850.n2 a_1129_n5850.n1 4.517
R21878 a_7067_n1053.t0 a_7067_n1053.t1 242.857
R21879 Din[2].n0 Din[2].t0 215.292
R21880 Din[2].n0 Din[2].t1 187.376
R21881 Din[2] Din[2].n0 84.902
R21882 a_5917_4148.t0 a_5917_4148.t1 242.857
R21883 a_11846_n7203.n0 a_11846_n7203.t1 63.08
R21884 a_11846_n7203.t0 a_11846_n7203.n0 41.306
R21885 a_11846_n7203.n0 a_11846_n7203.t2 2.251
R21886 a_11984_n7203.t0 a_11984_n7203.t1 68.741
R21887 a_5193_n2086.t0 a_5193_n2086.t1 34.8
R21888 a_2015_1698.t0 a_2015_1698.t1 242.857
R21889 a_4890_2662.t0 a_4890_2662.t1 242.857
R21890 a_7190_3184.t0 a_7190_3184.t1 242.857
R21891 a_742_n30.t0 a_742_n30.t1 242.857
R21892 a_5527_n2234.n2 a_5527_n2234.t0 282.97
R21893 a_5527_n2234.n1 a_5527_n2234.t4 240.683
R21894 a_5527_n2234.n0 a_5527_n2234.t2 209.208
R21895 a_5527_n2234.n0 a_5527_n2234.t3 194.167
R21896 a_5527_n2234.t1 a_5527_n2234.n2 183.404
R21897 a_5527_n2234.n1 a_5527_n2234.n0 14.805
R21898 a_5527_n2234.n2 a_5527_n2234.n1 6.415
R21899 a_5650_n2132.n0 a_5650_n2132.t2 489.336
R21900 a_5650_n2132.n0 a_5650_n2132.t1 243.258
R21901 a_5650_n2132.t0 a_5650_n2132.n0 214.415
R21902 a_n1495_n6849.t0 a_n1495_n6849.t1 42.707
R21903 a_n1460_n6503.n0 a_n1460_n6503.t0 65.064
R21904 a_n1460_n6503.n0 a_n1460_n6503.t2 42.011
R21905 a_n1460_n6503.t1 a_n1460_n6503.n0 2.113
R21906 ADC7_OUT[1].n0 ADC7_OUT[1].t4 1355.37
R21907 ADC7_OUT[1].n0 ADC7_OUT[1].t3 820.859
R21908 ADC7_OUT[1].n3 ADC7_OUT[1].t0 338.173
R21909 ADC7_OUT[1].n2 ADC7_OUT[1].t1 266.644
R21910 ADC7_OUT[1].n1 ADC7_OUT[1].n0 149.035
R21911 ADC7_OUT[1] ADC7_OUT[1].n3 45.977
R21912 ADC7_OUT[1].n1 ADC7_OUT[1].t2 45.968
R21913 ADC7_OUT[1].n3 ADC7_OUT[1].n2 45.929
R21914 ADC7_OUT[1].n2 ADC7_OUT[1].n1 17.317
R21915 a_290_2421.t0 a_290_2421.t1 242.857
R21916 a_n2148_n4114.t1 a_n2148_n4114.t0 336.812
R21917 a_n2207_n4470.t0 a_n2207_n4470.t1 68.741
R21918 Din[7].n0 Din[7].t0 215.292
R21919 Din[7].n0 Din[7].t1 187.376
R21920 Din[7] Din[7].n0 84.876
R21921 a_290_n271.t0 a_290_n271.t1 242.857
R21922 a_4192_2421.t0 a_4192_2421.t1 242.857
R21923 a_11549_n8026.n0 a_11549_n8026.t0 65.063
R21924 a_11549_n8026.n0 a_11549_n8026.t2 42.011
R21925 a_11549_n8026.t1 a_11549_n8026.n0 2.113
R21926 a_4192_n271.t0 a_4192_n271.t1 242.857
R21927 a_5465_2421.t0 a_5465_2421.t1 242.857
R21928 a_8327_2406.n0 a_8327_2406.t1 362.857
R21929 a_8327_2406.t5 a_8327_2406.t3 337.399
R21930 a_8327_2406.t3 a_8327_2406.t4 298.839
R21931 a_8327_2406.n0 a_8327_2406.t5 280.405
R21932 a_8327_2406.n1 a_8327_2406.t2 200
R21933 a_8327_2406.n1 a_8327_2406.n0 172.311
R21934 a_8327_2406.n2 a_8327_2406.n1 24
R21935 a_8327_2406.n1 a_8327_2406.t0 21.212
R21936 a_1440_1457.t0 a_1440_1457.t1 242.857
R21937 a_13033_n5338.n0 a_13033_n5338.t0 63.08
R21938 a_13033_n5338.n0 a_13033_n5338.t2 41.307
R21939 a_13033_n5338.t1 a_13033_n5338.n0 2.251
R21940 a_3822_3184.n0 a_3822_3184.t1 358.166
R21941 a_3822_3184.t4 a_3822_3184.t3 337.399
R21942 a_3822_3184.t3 a_3822_3184.t5 285.986
R21943 a_3822_3184.n0 a_3822_3184.t4 282.573
R21944 a_3822_3184.n1 a_3822_3184.t0 202.857
R21945 a_3822_3184.n1 a_3822_3184.n0 173.817
R21946 a_3822_3184.n1 a_3822_3184.t2 20.826
R21947 a_3822_3184.n2 a_3822_3184.n1 20.689
R21948 a_3727_3169.n0 a_3727_3169.t2 362.857
R21949 a_3727_3169.t3 a_3727_3169.t4 337.399
R21950 a_3727_3169.t4 a_3727_3169.t5 298.839
R21951 a_3727_3169.n0 a_3727_3169.t3 280.405
R21952 a_3727_3169.n1 a_3727_3169.t0 200
R21953 a_3727_3169.n1 a_3727_3169.n0 172.311
R21954 a_3727_3169.n2 a_3727_3169.n1 24
R21955 a_3727_3169.n1 a_3727_3169.t1 21.212
R21956 RWLB[4].n0 RWLB[4].t3 154.228
R21957 RWLB[4].n14 RWLB[4].t4 149.249
R21958 RWLB[4].n13 RWLB[4].t6 149.249
R21959 RWLB[4].n12 RWLB[4].t1 149.249
R21960 RWLB[4].n11 RWLB[4].t11 149.249
R21961 RWLB[4].n10 RWLB[4].t5 149.249
R21962 RWLB[4].n9 RWLB[4].t8 149.249
R21963 RWLB[4].n8 RWLB[4].t9 149.249
R21964 RWLB[4].n7 RWLB[4].t14 149.249
R21965 RWLB[4].n6 RWLB[4].t7 149.249
R21966 RWLB[4].n5 RWLB[4].t12 149.249
R21967 RWLB[4].n4 RWLB[4].t13 149.249
R21968 RWLB[4].n3 RWLB[4].t2 149.249
R21969 RWLB[4].n2 RWLB[4].t10 149.249
R21970 RWLB[4].n1 RWLB[4].t0 149.249
R21971 RWLB[4].n0 RWLB[4].t15 149.249
R21972 RWLB[4] RWLB[4].n14 47.816
R21973 RWLB[4].n1 RWLB[4].n0 4.979
R21974 RWLB[4].n2 RWLB[4].n1 4.979
R21975 RWLB[4].n3 RWLB[4].n2 4.979
R21976 RWLB[4].n4 RWLB[4].n3 4.979
R21977 RWLB[4].n5 RWLB[4].n4 4.979
R21978 RWLB[4].n6 RWLB[4].n5 4.979
R21979 RWLB[4].n7 RWLB[4].n6 4.979
R21980 RWLB[4].n8 RWLB[4].n7 4.979
R21981 RWLB[4].n9 RWLB[4].n8 4.979
R21982 RWLB[4].n10 RWLB[4].n9 4.979
R21983 RWLB[4].n11 RWLB[4].n10 4.979
R21984 RWLB[4].n12 RWLB[4].n11 4.979
R21985 RWLB[4].n13 RWLB[4].n12 4.979
R21986 RWLB[4].n14 RWLB[4].n13 4.979
R21987 a_8217_2662.t0 a_8217_2662.t1 242.857
R21988 a_8327_n286.n0 a_8327_n286.t0 362.857
R21989 a_8327_n286.t5 a_8327_n286.t3 337.399
R21990 a_8327_n286.t3 a_8327_n286.t4 298.839
R21991 a_8327_n286.n0 a_8327_n286.t5 280.405
R21992 a_8327_n286.n1 a_8327_n286.t1 200
R21993 a_8327_n286.n1 a_8327_n286.n0 172.311
R21994 a_8327_n286.n2 a_8327_n286.n1 24
R21995 a_8327_n286.n1 a_8327_n286.t2 21.212
R21996 a_8422_n271.n0 a_8422_n271.t1 358.166
R21997 a_8422_n271.t3 a_8422_n271.t5 337.399
R21998 a_8422_n271.t5 a_8422_n271.t4 285.986
R21999 a_8422_n271.n0 a_8422_n271.t3 282.573
R22000 a_8422_n271.n1 a_8422_n271.t2 202.857
R22001 a_8422_n271.n1 a_8422_n271.n0 173.817
R22002 a_8422_n271.n1 a_8422_n271.t0 20.826
R22003 a_8422_n271.n2 a_8422_n271.n1 20.689
R22004 a_8902_n286.n0 a_8902_n286.t2 362.857
R22005 a_8902_n286.t5 a_8902_n286.t4 337.399
R22006 a_8902_n286.t4 a_8902_n286.t3 298.839
R22007 a_8902_n286.n0 a_8902_n286.t5 280.405
R22008 a_8902_n286.n1 a_8902_n286.t0 200
R22009 a_8902_n286.n1 a_8902_n286.n0 172.311
R22010 a_8902_n286.n2 a_8902_n286.n1 24
R22011 a_8902_n286.n1 a_8902_n286.t1 21.212
R22012 a_6122_4686.n0 a_6122_4686.t1 358.166
R22013 a_6122_4686.t3 a_6122_4686.t5 337.399
R22014 a_6122_4686.t5 a_6122_4686.t4 285.986
R22015 a_6122_4686.n0 a_6122_4686.t3 282.573
R22016 a_6122_4686.n1 a_6122_4686.t2 202.857
R22017 a_6122_4686.n1 a_6122_4686.n0 173.817
R22018 a_6122_4686.n1 a_6122_4686.t0 20.826
R22019 a_6122_4686.n2 a_6122_4686.n1 20.689
R22020 ADC2_OUT[1].n0 ADC2_OUT[1].t4 1355.37
R22021 ADC2_OUT[1].n0 ADC2_OUT[1].t3 820.859
R22022 ADC2_OUT[1].n3 ADC2_OUT[1].t0 335.914
R22023 ADC2_OUT[1].n2 ADC2_OUT[1].t1 266.644
R22024 ADC2_OUT[1].n1 ADC2_OUT[1].n0 149.035
R22025 ADC2_OUT[1].n3 ADC2_OUT[1].n2 48.188
R22026 ADC2_OUT[1].n1 ADC2_OUT[1].t2 45.968
R22027 ADC2_OUT[1] ADC2_OUT[1].n3 45.633
R22028 ADC2_OUT[1].n2 ADC2_OUT[1].n1 17.317
R22029 a_8525_n2132.n0 a_8525_n2132.t2 489.336
R22030 a_8525_n2132.n0 a_8525_n2132.t1 243.258
R22031 a_8525_n2132.t0 a_8525_n2132.n0 214.415
R22032 Din[4].n0 Din[4].t0 215.292
R22033 Din[4].n0 Din[4].t1 187.376
R22034 Din[4] Din[4].n0 84.903
R22035 a_8217_n1053.t0 a_8217_n1053.t1 242.857
R22036 a_6492_4148.t0 a_6492_4148.t1 242.857
R22037 a_6602_3169.n0 a_6602_3169.t1 362.857
R22038 a_6602_3169.t3 a_6602_3169.t5 337.399
R22039 a_6602_3169.t5 a_6602_3169.t4 298.839
R22040 a_6602_3169.n0 a_6602_3169.t3 280.405
R22041 a_6602_3169.n1 a_6602_3169.t0 200
R22042 a_6602_3169.n1 a_6602_3169.n0 172.311
R22043 a_6602_3169.n2 a_6602_3169.n1 24
R22044 a_6602_3169.n1 a_6602_3169.t2 21.212
R22045 a_8915_211.t0 a_8915_211.t1 242.857
R22046 a_7765_4148.t0 a_7765_4148.t1 242.857
R22047 a_1427_3892.n0 a_1427_3892.t2 362.857
R22048 a_1427_3892.t5 a_1427_3892.t3 337.399
R22049 a_1427_3892.t3 a_1427_3892.t4 298.839
R22050 a_1427_3892.n0 a_1427_3892.t5 280.405
R22051 a_1427_3892.n1 a_1427_3892.t0 200
R22052 a_1427_3892.n1 a_1427_3892.n0 172.311
R22053 a_1427_3892.n2 a_1427_3892.n1 24
R22054 a_1427_3892.n1 a_1427_3892.t1 21.212
R22055 a_2015_1216.t0 a_2015_1216.t1 242.857
R22056 a_2002_196.n0 a_2002_196.t2 362.857
R22057 a_2002_196.t3 a_2002_196.t5 337.399
R22058 a_2002_196.t5 a_2002_196.t4 298.839
R22059 a_2002_196.n0 a_2002_196.t3 280.405
R22060 a_2002_196.n1 a_2002_196.t0 200
R22061 a_2002_196.n1 a_2002_196.n0 172.311
R22062 a_2002_196.n2 a_2002_196.n1 24
R22063 a_2002_196.n1 a_2002_196.t1 21.212
R22064 a_2097_211.n0 a_2097_211.t1 358.166
R22065 a_2097_211.t4 a_2097_211.t3 337.399
R22066 a_2097_211.t3 a_2097_211.t5 285.986
R22067 a_2097_211.n0 a_2097_211.t4 282.573
R22068 a_2097_211.n1 a_2097_211.t2 202.857
R22069 a_2097_211.n1 a_2097_211.n0 173.817
R22070 a_2097_211.n1 a_2097_211.t0 20.826
R22071 a_2097_211.n2 a_2097_211.n1 20.689
R22072 a_2672_3184.n0 a_2672_3184.t1 358.166
R22073 a_2672_3184.t3 a_2672_3184.t4 337.399
R22074 a_2672_3184.t4 a_2672_3184.t5 285.986
R22075 a_2672_3184.n0 a_2672_3184.t3 282.573
R22076 a_2672_3184.n1 a_2672_3184.t0 202.857
R22077 a_2672_3184.n1 a_2672_3184.n0 173.817
R22078 a_2672_3184.n1 a_2672_3184.t2 20.826
R22079 a_2672_3184.n2 a_2672_3184.n1 20.689
R22080 a_2577_3169.n0 a_2577_3169.t2 362.857
R22081 a_2577_3169.t3 a_2577_3169.t4 337.399
R22082 a_2577_3169.t4 a_2577_3169.t5 298.839
R22083 a_2577_3169.n0 a_2577_3169.t3 280.405
R22084 a_2577_3169.n1 a_2577_3169.t0 200
R22085 a_2577_3169.n1 a_2577_3169.n0 172.311
R22086 a_2577_3169.n2 a_2577_3169.n1 24
R22087 a_2577_3169.n1 a_2577_3169.t1 21.212
R22088 a_3822_2943.n0 a_3822_2943.t2 358.166
R22089 a_3822_2943.t5 a_3822_2943.t4 337.399
R22090 a_3822_2943.t4 a_3822_2943.t3 285.986
R22091 a_3822_2943.n0 a_3822_2943.t5 282.573
R22092 a_3822_2943.n1 a_3822_2943.t0 202.857
R22093 a_3822_2943.n1 a_3822_2943.n0 173.817
R22094 a_3822_2943.n1 a_3822_2943.t1 20.826
R22095 a_3822_2943.n2 a_3822_2943.n1 20.689
R22096 a_9367_n812.t0 a_9367_n812.t1 242.857
R22097 a_7642_2421.t0 a_7642_2421.t1 242.857
R22098 a_7177_960.n0 a_7177_960.t2 362.857
R22099 a_7177_960.t3 a_7177_960.t5 337.399
R22100 a_7177_960.t5 a_7177_960.t4 298.839
R22101 a_7177_960.n0 a_7177_960.t3 280.405
R22102 a_7177_960.n1 a_7177_960.t0 200
R22103 a_7177_960.n1 a_7177_960.n0 172.311
R22104 a_7177_960.n2 a_7177_960.n1 24
R22105 a_7177_960.n1 a_7177_960.t1 21.212
R22106 a_1892_2180.t0 a_1892_2180.t1 242.857
R22107 a_7765_693.t0 a_7765_693.t1 242.857
R22108 a_1427_2406.n0 a_1427_2406.t2 362.857
R22109 a_1427_2406.t3 a_1427_2406.t4 337.399
R22110 a_1427_2406.t4 a_1427_2406.t5 298.839
R22111 a_1427_2406.n0 a_1427_2406.t3 280.405
R22112 a_1427_2406.n1 a_1427_2406.t0 200
R22113 a_1427_2406.n1 a_1427_2406.n0 172.311
R22114 a_1427_2406.n2 a_1427_2406.n1 24
R22115 a_1427_2406.n1 a_1427_2406.t1 21.212
R22116 a_7642_n271.t0 a_7642_n271.t1 242.857
R22117 a_7785_n1371.n1 a_7785_n1371.t4 550.94
R22118 a_7785_n1371.n1 a_7785_n1371.t3 500.621
R22119 a_7785_n1371.t2 a_7785_n1371.n2 192.787
R22120 a_7785_n1371.n0 a_7785_n1371.t0 163.997
R22121 a_7785_n1371.n2 a_7785_n1371.n1 149.035
R22122 a_7785_n1371.n0 a_7785_n1371.t1 54.068
R22123 a_7785_n1371.n2 a_7785_n1371.n0 17.317
R22124 SA_OUT[13].n1 SA_OUT[13].t4 661.027
R22125 SA_OUT[13].n1 SA_OUT[13].t3 392.255
R22126 SA_OUT[13].n2 SA_OUT[13].t2 223.716
R22127 SA_OUT[13].n0 SA_OUT[13].t0 153.977
R22128 SA_OUT[13].n2 SA_OUT[13].n1 143.764
R22129 SA_OUT[13].n0 SA_OUT[13].t1 59.86
R22130 SA_OUT[13] SA_OUT[13].n3 13.483
R22131 SA_OUT[13].n3 SA_OUT[13].n0 3.764
R22132 SA_OUT[13].n3 SA_OUT[13].n2 0.752
R22133 a_7765_3907.t0 a_7765_3907.t1 242.857
R22134 a_8915_2421.t0 a_8915_2421.t1 242.857
R22135 a_1427_n286.n0 a_1427_n286.t2 362.857
R22136 a_1427_n286.t3 a_1427_n286.t4 337.399
R22137 a_1427_n286.t4 a_1427_n286.t5 298.839
R22138 a_1427_n286.n0 a_1427_n286.t3 280.405
R22139 a_1427_n286.n1 a_1427_n286.t0 200
R22140 a_1427_n286.n1 a_1427_n286.n0 172.311
R22141 a_1427_n286.n2 a_1427_n286.n1 24
R22142 a_1427_n286.n1 a_1427_n286.t1 21.212
R22143 Din[9].n0 Din[9].t0 215.292
R22144 Din[9].n0 Din[9].t1 187.376
R22145 Din[9] Din[9].n0 84.894
R22146 a_6040_1939.t0 a_6040_1939.t1 242.857
R22147 a_4890_1939.t0 a_4890_1939.t1 242.857
R22148 a_8422_211.n0 a_8422_211.t1 358.166
R22149 a_8422_211.t4 a_8422_211.t3 337.399
R22150 a_8422_211.t3 a_8422_211.t5 285.986
R22151 a_8422_211.n0 a_8422_211.t4 282.573
R22152 a_8422_211.n1 a_8422_211.t0 202.857
R22153 a_8422_211.n1 a_8422_211.n0 173.817
R22154 a_8422_211.n1 a_8422_211.t2 20.826
R22155 a_8422_211.n2 a_8422_211.n1 20.689
R22156 a_8327_196.n0 a_8327_196.t2 362.857
R22157 a_8327_196.t3 a_8327_196.t5 337.399
R22158 a_8327_196.t5 a_8327_196.t4 298.839
R22159 a_8327_196.n0 a_8327_196.t3 280.405
R22160 a_8327_196.n1 a_8327_196.t0 200
R22161 a_8327_196.n1 a_8327_196.n0 172.311
R22162 a_8327_196.n2 a_8327_196.n1 24
R22163 a_8327_196.n1 a_8327_196.t1 21.212
R22164 a_947_n512.n0 a_947_n512.t2 358.166
R22165 a_947_n512.t4 a_947_n512.t5 337.399
R22166 a_947_n512.t5 a_947_n512.t3 285.986
R22167 a_947_n512.n0 a_947_n512.t4 282.573
R22168 a_947_n512.n1 a_947_n512.t0 202.857
R22169 a_947_n512.n1 a_947_n512.n0 173.817
R22170 a_947_n512.n1 a_947_n512.t1 20.826
R22171 a_947_n512.n2 a_947_n512.n1 20.689
R22172 a_2097_1939.n0 a_2097_1939.t1 358.166
R22173 a_2097_1939.t4 a_2097_1939.t5 337.399
R22174 a_2097_1939.t5 a_2097_1939.t3 285.986
R22175 a_2097_1939.n0 a_2097_1939.t4 282.573
R22176 a_2097_1939.n1 a_2097_1939.t2 202.857
R22177 a_2097_1939.n1 a_2097_1939.n0 173.817
R22178 a_2097_1939.n1 a_2097_1939.t0 20.826
R22179 a_2097_1939.n2 a_2097_1939.n1 20.689
R22180 a_2467_1939.t0 a_2467_1939.t1 242.857
R22181 a_8568_n2426.n3 a_8568_n2426.t3 475.39
R22182 a_8568_n2426.t5 a_8568_n2426.t7 228.696
R22183 a_8568_n2426.n3 a_8568_n2426.n2 198.34
R22184 a_8568_n2426.n2 a_8568_n2426.t1 185.704
R22185 a_8568_n2426.n0 a_8568_n2426.t5 126.761
R22186 a_8568_n2426.n1 a_8568_n2426.t6 126.284
R22187 a_8568_n2426.n1 a_8568_n2426.t0 126.284
R22188 a_8568_n2426.t2 a_8568_n2426.n3 124.375
R22189 a_8568_n2426.t0 a_8568_n2426.n0 115.122
R22190 a_8568_n2426.n0 a_8568_n2426.t4 111.229
R22191 a_8568_n2426.n2 a_8568_n2426.n1 8.764
R22192 a_12701_n5092.t0 a_12701_n5092.t1 42.705
R22193 a_5547_2421.n0 a_5547_2421.t0 358.166
R22194 a_5547_2421.t5 a_5547_2421.t3 337.399
R22195 a_5547_2421.t3 a_5547_2421.t4 285.986
R22196 a_5547_2421.n0 a_5547_2421.t5 282.573
R22197 a_5547_2421.n1 a_5547_2421.t2 202.857
R22198 a_5547_2421.n1 a_5547_2421.n0 173.817
R22199 a_5547_2421.n1 a_5547_2421.t1 20.826
R22200 a_5547_2421.n2 a_5547_2421.n1 20.689
R22201 a_5452_2406.n0 a_5452_2406.t2 362.857
R22202 a_5452_2406.t3 a_5452_2406.t4 337.399
R22203 a_5452_2406.t4 a_5452_2406.t5 298.839
R22204 a_5452_2406.n0 a_5452_2406.t3 280.405
R22205 a_5452_2406.n1 a_5452_2406.t0 200
R22206 a_5452_2406.n1 a_5452_2406.n0 172.311
R22207 a_5452_2406.n2 a_5452_2406.n1 24
R22208 a_5452_2406.n1 a_5452_2406.t1 21.212
R22209 a_6040_1698.t0 a_6040_1698.t1 242.857
R22210 a_11549_n5293.n0 a_11549_n5293.t0 65.063
R22211 a_11549_n5293.n0 a_11549_n5293.t2 42.011
R22212 a_11549_n5293.t1 a_11549_n5293.n0 2.113
R22213 ADC7_OUT[0].n0 ADC7_OUT[0].t3 1354.27
R22214 ADC7_OUT[0].n0 ADC7_OUT[0].t4 821.954
R22215 ADC7_OUT[0].n3 ADC7_OUT[0].t0 344.126
R22216 ADC7_OUT[0].n2 ADC7_OUT[0].t2 266.575
R22217 ADC7_OUT[0].n1 ADC7_OUT[0].n0 149.035
R22218 ADC7_OUT[0] ADC7_OUT[0].n3 61.829
R22219 ADC7_OUT[0].n1 ADC7_OUT[0].t1 46.723
R22220 ADC7_OUT[0].n3 ADC7_OUT[0].n2 39.905
R22221 ADC7_OUT[0].n2 ADC7_OUT[0].n1 17.317
R22222 a_4745_n4470.n0 a_4745_n4470.t1 63.08
R22223 a_4745_n4470.t0 a_4745_n4470.n0 41.306
R22224 a_4745_n4470.n0 a_4745_n4470.t2 2.251
R22225 a_4675_n4483.n0 a_4675_n4483.t3 1464.36
R22226 a_4675_n4483.n0 a_4675_n4483.t4 713.588
R22227 a_4675_n4483.n1 a_4675_n4483.t2 374.998
R22228 a_4675_n4483.n1 a_4675_n4483.t1 273.351
R22229 a_4675_n4483.n2 a_4675_n4483.n0 143.764
R22230 a_4675_n4483.t0 a_4675_n4483.n2 78.209
R22231 a_4675_n4483.n2 a_4675_n4483.n1 4.517
R22232 a_18_n4470.n0 a_18_n4470.t0 63.08
R22233 a_18_n4470.n0 a_18_n4470.t2 41.305
R22234 a_18_n4470.t1 a_18_n4470.n0 2.251
R22235 a_1427_3410.n0 a_1427_3410.t2 362.857
R22236 a_1427_3410.t5 a_1427_3410.t3 337.399
R22237 a_1427_3410.t3 a_1427_3410.t4 298.839
R22238 a_1427_3410.n0 a_1427_3410.t5 280.405
R22239 a_1427_3410.n1 a_1427_3410.t0 200
R22240 a_1427_3410.n1 a_1427_3410.n0 172.311
R22241 a_1427_3410.n2 a_1427_3410.n1 24
R22242 a_1427_3410.n1 a_1427_3410.t1 21.212
R22243 a_3042_2662.t0 a_3042_2662.t1 242.857
R22244 a_2467_1698.t0 a_2467_1698.t1 242.857
R22245 a_1317_3666.t0 a_1317_3666.t1 242.857
R22246 a_1440_4686.t0 a_1440_4686.t1 242.857
R22247 a_7067_211.t0 a_7067_211.t1 242.857
R22248 ADC13_OUT[3].n0 ADC13_OUT[3].t4 1355.37
R22249 ADC13_OUT[3].n0 ADC13_OUT[3].t3 820.859
R22250 ADC13_OUT[3].n3 ADC13_OUT[3].t0 327.632
R22251 ADC13_OUT[3].n2 ADC13_OUT[3].t1 266.644
R22252 ADC13_OUT[3].n1 ADC13_OUT[3].n0 149.035
R22253 ADC13_OUT[3].n3 ADC13_OUT[3].n2 56.47
R22254 ADC13_OUT[3].n1 ADC13_OUT[3].t2 45.968
R22255 ADC13_OUT[3] ADC13_OUT[3].n3 22.356
R22256 ADC13_OUT[3].n2 ADC13_OUT[3].n1 17.317
R22257 a_11776_n8583.n0 a_11776_n8583.t4 1465.51
R22258 a_11776_n8583.n0 a_11776_n8583.t3 712.44
R22259 a_11776_n8583.n1 a_11776_n8583.t0 375.067
R22260 a_11776_n8583.n1 a_11776_n8583.t2 272.668
R22261 a_11776_n8583.n2 a_11776_n8583.n0 143.764
R22262 a_11776_n8583.t1 a_11776_n8583.n2 78.193
R22263 a_11776_n8583.n2 a_11776_n8583.n1 4.517
R22264 EN.n13 EN.t5 318.889
R22265 EN.n14 EN.t10 317.428
R22266 EN.n11 EN.t11 315.125
R22267 EN.n12 EN.t3 313.664
R22268 EN.n7 EN.t6 310.446
R22269 EN.n3 EN.t0 310.058
R22270 EN.n0 EN.t13 309.917
R22271 EN.n1 EN.t1 308.919
R22272 EN.n5 EN.t7 308.919
R22273 EN.n9 EN.t12 308.919
R22274 EN.n8 EN.t14 308.621
R22275 EN.n4 EN.t8 308.21
R22276 EN.n2 EN.t9 307.845
R22277 EN.n6 EN.t15 307.845
R22278 EN.n10 EN.t4 307.458
R22279 EN.n0 EN.t2 306.705
R22280 EN EN.n14 8.279
R22281 EN.n3 EN.n2 1.549
R22282 EN.n1 EN.n0 1.546
R22283 EN.n5 EN.n4 1.546
R22284 EN.n11 EN.n10 1.545
R22285 EN.n13 EN.n12 1.545
R22286 EN.n7 EN.n6 1.542
R22287 EN.n9 EN.n8 1.542
R22288 EN.n8 EN.n7 0.235
R22289 EN.n6 EN.n5 0.229
R22290 EN.n12 EN.n11 0.229
R22291 EN.n14 EN.n13 0.229
R22292 EN.n10 EN.n9 0.227
R22293 EN.n2 EN.n1 0.226
R22294 EN.n4 EN.n3 0.226
R22295 a_7765_3425.t0 a_7765_3425.t1 242.857
R22296 a_8902_960.n0 a_8902_960.t1 362.857
R22297 a_8902_960.t3 a_8902_960.t5 337.399
R22298 a_8902_960.t5 a_8902_960.t4 298.839
R22299 a_8902_960.n0 a_8902_960.t3 280.405
R22300 a_8902_960.n1 a_8902_960.t0 200
R22301 a_8902_960.n1 a_8902_960.n0 172.311
R22302 a_8902_960.n2 a_8902_960.n1 24
R22303 a_8902_960.n1 a_8902_960.t2 21.212
R22304 a_8997_975.n0 a_8997_975.t1 358.166
R22305 a_8997_975.t4 a_8997_975.t5 337.399
R22306 a_8997_975.t5 a_8997_975.t3 285.986
R22307 a_8997_975.n0 a_8997_975.t4 282.573
R22308 a_8997_975.n1 a_8997_975.t2 202.857
R22309 a_8997_975.n1 a_8997_975.n0 173.817
R22310 a_8997_975.n1 a_8997_975.t0 20.826
R22311 a_8997_975.n2 a_8997_975.n1 20.689
R22312 SA_OUT[15].n1 SA_OUT[15].t4 661.027
R22313 SA_OUT[15].n1 SA_OUT[15].t3 392.255
R22314 SA_OUT[15].n2 SA_OUT[15].t0 223.716
R22315 SA_OUT[15].n0 SA_OUT[15].t2 153.977
R22316 SA_OUT[15].n2 SA_OUT[15].n1 143.764
R22317 SA_OUT[15].n0 SA_OUT[15].t1 59.86
R22318 SA_OUT[15] SA_OUT[15].n3 13.188
R22319 SA_OUT[15].n3 SA_OUT[15].n2 3.011
R22320 SA_OUT[15].n3 SA_OUT[15].n0 1.505
R22321 a_1522_2421.n0 a_1522_2421.t2 358.166
R22322 a_1522_2421.t3 a_1522_2421.t5 337.399
R22323 a_1522_2421.t5 a_1522_2421.t4 285.986
R22324 a_1522_2421.n0 a_1522_2421.t3 282.573
R22325 a_1522_2421.n1 a_1522_2421.t0 202.857
R22326 a_1522_2421.n1 a_1522_2421.n0 173.817
R22327 a_1522_2421.n1 a_1522_2421.t1 20.826
R22328 a_1522_2421.n2 a_1522_2421.n1 20.689
R22329 a_9405_n5850.n0 a_9405_n5850.t4 1465.51
R22330 a_9405_n5850.n0 a_9405_n5850.t3 712.44
R22331 a_9405_n5850.n1 a_9405_n5850.t0 375.067
R22332 a_9405_n5850.n1 a_9405_n5850.t1 272.668
R22333 a_9405_n5850.n2 a_9405_n5850.n0 143.764
R22334 a_9405_n5850.t2 a_9405_n5850.n2 78.193
R22335 a_9405_n5850.n2 a_9405_n5850.n1 4.517
R22336 a_11846_n4470.n0 a_11846_n4470.t0 63.08
R22337 a_11846_n4470.t1 a_11846_n4470.n0 41.306
R22338 a_11846_n4470.n0 a_11846_n4470.t2 2.251
R22339 a_11984_n4470.t0 a_11984_n4470.t1 68.741
R22340 a_6027_2647.n0 a_6027_2647.t0 362.857
R22341 a_6027_2647.t3 a_6027_2647.t4 337.399
R22342 a_6027_2647.t4 a_6027_2647.t5 298.839
R22343 a_6027_2647.n0 a_6027_2647.t3 280.405
R22344 a_6027_2647.n1 a_6027_2647.t2 200
R22345 a_6027_2647.n1 a_6027_2647.n0 172.311
R22346 a_6027_2647.n2 a_6027_2647.n1 24
R22347 a_6027_2647.n1 a_6027_2647.t1 21.212
R22348 a_5547_1939.n0 a_5547_1939.t1 358.166
R22349 a_5547_1939.t4 a_5547_1939.t5 337.399
R22350 a_5547_1939.t5 a_5547_1939.t3 285.986
R22351 a_5547_1939.n0 a_5547_1939.t4 282.573
R22352 a_5547_1939.n1 a_5547_1939.t2 202.857
R22353 a_5547_1939.n1 a_5547_1939.n0 173.817
R22354 a_5547_1939.n1 a_5547_1939.t0 20.826
R22355 a_5547_1939.n2 a_5547_1939.n1 20.689
R22356 a_5917_1939.t0 a_5917_1939.t1 242.857
R22357 a_8792_211.t0 a_8792_211.t1 242.857
R22358 a_n1233_n8583.n0 a_n1233_n8583.t4 1465.51
R22359 a_n1233_n8583.n0 a_n1233_n8583.t3 712.44
R22360 a_n1233_n8583.n1 a_n1233_n8583.t0 375.067
R22361 a_n1233_n8583.n1 a_n1233_n8583.t1 272.668
R22362 a_n1233_n8583.n2 a_n1233_n8583.n0 143.764
R22363 a_n1233_n8583.t2 a_n1233_n8583.n2 78.193
R22364 a_n1233_n8583.n2 a_n1233_n8583.n1 4.517
R22365 a_n3565_n4483.n0 a_n3565_n4483.t3 1464.36
R22366 a_n3565_n4483.n0 a_n3565_n4483.t4 713.588
R22367 a_n3565_n4483.n1 a_n3565_n4483.t0 374.998
R22368 a_n3565_n4483.n1 a_n3565_n4483.t2 273.351
R22369 a_n3565_n4483.n2 a_n3565_n4483.n0 143.764
R22370 a_n3565_n4483.t1 a_n3565_n4483.n2 78.209
R22371 a_n3565_n4483.n2 a_n3565_n4483.n1 4.517
R22372 ADC0_OUT[0].n0 ADC0_OUT[0].t3 1354.27
R22373 ADC0_OUT[0].n0 ADC0_OUT[0].t4 821.954
R22374 ADC0_OUT[0].n3 ADC0_OUT[0].t0 334.338
R22375 ADC0_OUT[0].n2 ADC0_OUT[0].t1 266.575
R22376 ADC0_OUT[0].n1 ADC0_OUT[0].n0 149.035
R22377 ADC0_OUT[0] ADC0_OUT[0].n3 61.883
R22378 ADC0_OUT[0].n3 ADC0_OUT[0].n2 49.694
R22379 ADC0_OUT[0].n1 ADC0_OUT[0].t2 46.723
R22380 ADC0_OUT[0].n2 ADC0_OUT[0].n1 17.317
R22381 a_2015_4445.t0 a_2015_4445.t1 242.857
R22382 a_1892_1457.t0 a_1892_1457.t1 242.857
R22383 a_7272_693.n0 a_7272_693.t2 358.166
R22384 a_7272_693.t5 a_7272_693.t4 337.399
R22385 a_7272_693.t4 a_7272_693.t3 285.986
R22386 a_7272_693.n0 a_7272_693.t5 282.573
R22387 a_7272_693.n1 a_7272_693.t0 202.857
R22388 a_7272_693.n1 a_7272_693.n0 173.817
R22389 a_7272_693.n1 a_7272_693.t1 20.826
R22390 a_7272_693.n2 a_7272_693.n1 20.689
R22391 a_290_452.t0 a_290_452.t1 242.857
R22392 a_7835_n1770.n0 a_7835_n1770.t2 325.682
R22393 a_7835_n1770.n0 a_7835_n1770.t1 322.294
R22394 a_7835_n1770.t0 a_7835_n1770.n0 73.623
R22395 a_2590_3907.t0 a_2590_3907.t1 242.857
R22396 a_6040_1216.t0 a_6040_1216.t1 242.857
R22397 a_742_n512.t0 a_742_n512.t1 242.857
R22398 a_n1495_n4116.t0 a_n1495_n4116.t1 42.707
R22399 a_n1460_n3770.n0 a_n1460_n3770.t0 65.064
R22400 a_n1460_n3770.n0 a_n1460_n3770.t2 42.011
R22401 a_n1460_n3770.t1 a_n1460_n3770.n0 2.113
R22402 a_6697_3184.n0 a_6697_3184.t2 358.166
R22403 a_6697_3184.t3 a_6697_3184.t4 337.399
R22404 a_6697_3184.t4 a_6697_3184.t5 285.986
R22405 a_6697_3184.n0 a_6697_3184.t3 282.573
R22406 a_6697_3184.n1 a_6697_3184.t0 202.857
R22407 a_6697_3184.n1 a_6697_3184.n0 173.817
R22408 a_6697_3184.n1 a_6697_3184.t1 20.826
R22409 a_6697_3184.n2 a_6697_3184.n1 20.689
R22410 a_5917_1698.t0 a_5917_1698.t1 242.857
R22411 a_3042_975.t0 a_3042_975.t1 242.857
R22412 a_7067_2180.t0 a_7067_2180.t1 242.857
R22413 a_3165_211.t0 a_3165_211.t1 242.857
R22414 a_2467_1216.t0 a_2467_1216.t1 242.857
R22415 a_2577_960.n0 a_2577_960.t2 362.857
R22416 a_2577_960.t3 a_2577_960.t5 337.399
R22417 a_2577_960.t5 a_2577_960.t4 298.839
R22418 a_2577_960.n0 a_2577_960.t3 280.405
R22419 a_2577_960.n1 a_2577_960.t0 200
R22420 a_2577_960.n1 a_2577_960.n0 172.311
R22421 a_2577_960.n2 a_2577_960.n1 24
R22422 a_2577_960.n1 a_2577_960.t1 21.212
R22423 a_2672_975.n0 a_2672_975.t2 358.166
R22424 a_2672_975.t5 a_2672_975.t3 337.399
R22425 a_2672_975.t3 a_2672_975.t4 285.986
R22426 a_2672_975.n0 a_2672_975.t5 282.573
R22427 a_2672_975.n1 a_2672_975.t0 202.857
R22428 a_2672_975.n1 a_2672_975.n0 173.817
R22429 a_2672_975.n1 a_2672_975.t1 20.826
R22430 a_2672_975.n2 a_2672_975.n1 20.689
R22431 a_3740_n1053.t0 a_3740_n1053.t1 242.857
R22432 a_4315_452.t0 a_4315_452.t1 242.857
R22433 a_3165_3666.t0 a_3165_3666.t1 242.857
R22434 a_6027_3651.n0 a_6027_3651.t1 362.857
R22435 a_6027_3651.t5 a_6027_3651.t3 337.399
R22436 a_6027_3651.t3 a_6027_3651.t4 298.839
R22437 a_6027_3651.n0 a_6027_3651.t5 280.405
R22438 a_6027_3651.n1 a_6027_3651.t2 200
R22439 a_6027_3651.n1 a_6027_3651.n0 172.311
R22440 a_6027_3651.n2 a_6027_3651.n1 24
R22441 a_6027_3651.n1 a_6027_3651.t0 21.212
R22442 a_2311_n7216.n0 a_2311_n7216.t4 1464.36
R22443 a_2311_n7216.n0 a_2311_n7216.t3 713.588
R22444 a_2311_n7216.n1 a_2311_n7216.t0 374.998
R22445 a_2311_n7216.n1 a_2311_n7216.t1 273.351
R22446 a_2311_n7216.n2 a_2311_n7216.n0 143.764
R22447 a_2311_n7216.t2 a_2311_n7216.n2 78.209
R22448 a_2311_n7216.n2 a_2311_n7216.n1 4.517
R22449 ADC5_OUT[2].n0 ADC5_OUT[2].t4 1354.27
R22450 ADC5_OUT[2].n0 ADC5_OUT[2].t3 821.954
R22451 ADC5_OUT[2].n3 ADC5_OUT[2].t0 349.397
R22452 ADC5_OUT[2].n2 ADC5_OUT[2].t2 266.575
R22453 ADC5_OUT[2].n1 ADC5_OUT[2].n0 149.035
R22454 ADC5_OUT[2].n1 ADC5_OUT[2].t1 46.723
R22455 ADC5_OUT[2] ADC5_OUT[2].n3 37.869
R22456 ADC5_OUT[2].n3 ADC5_OUT[2].n2 34.635
R22457 ADC5_OUT[2].n2 ADC5_OUT[2].n1 17.317
R22458 a_7272_2943.n0 a_7272_2943.t1 358.166
R22459 a_7272_2943.t3 a_7272_2943.t5 337.399
R22460 a_7272_2943.t5 a_7272_2943.t4 285.986
R22461 a_7272_2943.n0 a_7272_2943.t3 282.573
R22462 a_7272_2943.n1 a_7272_2943.t0 202.857
R22463 a_7272_2943.n1 a_7272_2943.n0 173.817
R22464 a_7272_2943.n1 a_7272_2943.t2 20.826
R22465 a_7272_2943.n2 a_7272_2943.n1 20.689
R22466 a_7177_2928.n0 a_7177_2928.t2 362.857
R22467 a_7177_2928.t3 a_7177_2928.t4 337.399
R22468 a_7177_2928.t4 a_7177_2928.t5 298.839
R22469 a_7177_2928.n0 a_7177_2928.t3 280.405
R22470 a_7177_2928.n1 a_7177_2928.t0 200
R22471 a_7177_2928.n1 a_7177_2928.n0 172.311
R22472 a_7177_2928.n2 a_7177_2928.n1 24
R22473 a_7177_2928.n1 a_7177_2928.t1 21.212
R22474 a_4890_211.t0 a_4890_211.t1 242.857
R22475 RWLB[3].n0 RWLB[3].t3 154.228
R22476 RWLB[3].n14 RWLB[3].t4 149.249
R22477 RWLB[3].n13 RWLB[3].t6 149.249
R22478 RWLB[3].n12 RWLB[3].t1 149.249
R22479 RWLB[3].n11 RWLB[3].t11 149.249
R22480 RWLB[3].n10 RWLB[3].t5 149.249
R22481 RWLB[3].n9 RWLB[3].t8 149.249
R22482 RWLB[3].n8 RWLB[3].t9 149.249
R22483 RWLB[3].n7 RWLB[3].t14 149.249
R22484 RWLB[3].n6 RWLB[3].t7 149.249
R22485 RWLB[3].n5 RWLB[3].t12 149.249
R22486 RWLB[3].n4 RWLB[3].t13 149.249
R22487 RWLB[3].n3 RWLB[3].t2 149.249
R22488 RWLB[3].n2 RWLB[3].t10 149.249
R22489 RWLB[3].n1 RWLB[3].t0 149.249
R22490 RWLB[3].n0 RWLB[3].t15 149.249
R22491 RWLB[3] RWLB[3].n14 47.816
R22492 RWLB[3].n1 RWLB[3].n0 4.979
R22493 RWLB[3].n2 RWLB[3].n1 4.979
R22494 RWLB[3].n3 RWLB[3].n2 4.979
R22495 RWLB[3].n4 RWLB[3].n3 4.979
R22496 RWLB[3].n5 RWLB[3].n4 4.979
R22497 RWLB[3].n6 RWLB[3].n5 4.979
R22498 RWLB[3].n7 RWLB[3].n6 4.979
R22499 RWLB[3].n8 RWLB[3].n7 4.979
R22500 RWLB[3].n9 RWLB[3].n8 4.979
R22501 RWLB[3].n10 RWLB[3].n9 4.979
R22502 RWLB[3].n11 RWLB[3].n10 4.979
R22503 RWLB[3].n12 RWLB[3].n11 4.979
R22504 RWLB[3].n13 RWLB[3].n12 4.979
R22505 RWLB[3].n14 RWLB[3].n13 4.979
R22506 a_8217_2943.t0 a_8217_2943.t1 242.857
R22507 a_3042_1939.t0 a_3042_1939.t1 242.857
R22508 a_6492_1939.t0 a_6492_1939.t1 242.857
R22509 a_2590_n271.t0 a_2590_n271.t1 242.857
R22510 a_372_2943.n0 a_372_2943.t2 358.166
R22511 a_372_2943.t5 a_372_2943.t4 337.399
R22512 a_372_2943.t4 a_372_2943.t3 285.986
R22513 a_372_2943.n0 a_372_2943.t5 282.573
R22514 a_372_2943.n1 a_372_2943.t0 202.857
R22515 a_372_2943.n1 a_372_2943.n0 173.817
R22516 a_372_2943.n1 a_372_2943.t1 20.826
R22517 a_372_2943.n2 a_372_2943.n1 20.689
R22518 a_742_2943.t0 a_742_2943.t1 242.857
R22519 a_6122_2662.n0 a_6122_2662.t1 358.166
R22520 a_6122_2662.t3 a_6122_2662.t5 337.399
R22521 a_6122_2662.t5 a_6122_2662.t4 285.986
R22522 a_6122_2662.n0 a_6122_2662.t3 282.573
R22523 a_6122_2662.n1 a_6122_2662.t2 202.857
R22524 a_6122_2662.n1 a_6122_2662.n0 173.817
R22525 a_6122_2662.n1 a_6122_2662.t0 20.826
R22526 a_6122_2662.n2 a_6122_2662.n1 20.689
R22527 a_3740_975.t0 a_3740_975.t1 242.857
R22528 a_2590_3425.t0 a_2590_3425.t1 242.857
R22529 a_5342_3666.t0 a_5342_3666.t1 242.857
R22530 a_6492_1698.t0 a_6492_1698.t1 242.857
R22531 a_5917_1216.t0 a_5917_1216.t1 242.857
R22532 a_n966_n8026.t1 a_n966_n8026.t0 336.814
R22533 a_n1025_n8071.t0 a_n1025_n8071.t1 68.74
R22534 a_5630_n8026.n0 a_5630_n8026.t0 65.063
R22535 a_5630_n8026.n0 a_5630_n8026.t2 42.011
R22536 a_5630_n8026.t1 a_5630_n8026.n0 2.113
R22537 a_1317_n1053.t0 a_1317_n1053.t1 242.857
R22538 a_6615_3666.t0 a_6615_3666.t1 242.857
R22539 a_7765_1698.t0 a_7765_1698.t1 242.857
R22540 a_2467_211.t0 a_2467_211.t1 242.857
R22541 a_5547_452.n0 a_5547_452.t0 358.166
R22542 a_5547_452.t5 a_5547_452.t4 337.399
R22543 a_5547_452.t4 a_5547_452.t3 285.986
R22544 a_5547_452.n0 a_5547_452.t5 282.573
R22545 a_5547_452.n1 a_5547_452.t2 202.857
R22546 a_5547_452.n1 a_5547_452.n0 173.817
R22547 a_5547_452.n1 a_5547_452.t1 20.826
R22548 a_5547_452.n2 a_5547_452.n1 20.689
R22549 a_5917_452.t0 a_5917_452.t1 242.857
R22550 a_7994_n8026.n0 a_7994_n8026.t0 65.063
R22551 a_7994_n8026.n0 a_7994_n8026.t2 42.011
R22552 a_7994_n8026.t1 a_7994_n8026.n0 2.113
R22553 a_4302_960.n0 a_4302_960.t2 362.857
R22554 a_4302_960.t3 a_4302_960.t5 337.399
R22555 a_4302_960.t5 a_4302_960.t4 298.839
R22556 a_4302_960.n0 a_4302_960.t3 280.405
R22557 a_4302_960.n1 a_4302_960.t0 200
R22558 a_4302_960.n1 a_4302_960.n0 172.311
R22559 a_4302_960.n2 a_4302_960.n1 24
R22560 a_4302_960.n1 a_4302_960.t1 21.212
R22561 a_7765_n812.t0 a_7765_n812.t1 242.857
R22562 a_1892_4686.t0 a_1892_4686.t1 242.857
R22563 a_7067_1457.t0 a_7067_1457.t1 242.857
R22564 a_2578_n6847.t1 a_2578_n6847.t0 336.812
R22565 a_2381_n7203.n0 a_2381_n7203.t0 63.08
R22566 a_2381_n7203.n0 a_2381_n7203.t2 41.305
R22567 a_2381_n7203.t1 a_2381_n7203.n0 2.251
R22568 a_2672_2180.n0 a_2672_2180.t1 358.166
R22569 a_2672_2180.t5 a_2672_2180.t3 337.399
R22570 a_2672_2180.t3 a_2672_2180.t4 285.986
R22571 a_2672_2180.n0 a_2672_2180.t5 282.573
R22572 a_2672_2180.n1 a_2672_2180.t2 202.857
R22573 a_2672_2180.n1 a_2672_2180.n0 173.817
R22574 a_2672_2180.n1 a_2672_2180.t0 20.826
R22575 a_2672_2180.n2 a_2672_2180.n1 20.689
R22576 a_852_1442.n0 a_852_1442.t0 362.857
R22577 a_852_1442.t3 a_852_1442.t4 337.399
R22578 a_852_1442.t4 a_852_1442.t5 298.839
R22579 a_852_1442.n0 a_852_1442.t3 280.405
R22580 a_852_1442.n1 a_852_1442.t2 200
R22581 a_852_1442.n1 a_852_1442.n0 172.311
R22582 a_852_1442.n2 a_852_1442.n1 24
R22583 a_852_1442.n1 a_852_1442.t1 21.212
R22584 a_6040_4445.t0 a_6040_4445.t1 242.857
R22585 a_2672_693.n0 a_2672_693.t2 358.166
R22586 a_2672_693.t5 a_2672_693.t4 337.399
R22587 a_2672_693.t4 a_2672_693.t3 285.986
R22588 a_2672_693.n0 a_2672_693.t5 282.573
R22589 a_2672_693.n1 a_2672_693.t0 202.857
R22590 a_2672_693.n1 a_2672_693.n0 173.817
R22591 a_2672_693.n1 a_2672_693.t1 20.826
R22592 a_2672_693.n2 a_2672_693.n1 20.689
R22593 a_5465_n30.t0 a_5465_n30.t1 242.857
R22594 a_2467_4445.t0 a_2467_4445.t1 242.857
R22595 a_947_1457.n0 a_947_1457.t1 358.166
R22596 a_947_1457.t4 a_947_1457.t5 337.399
R22597 a_947_1457.t5 a_947_1457.t3 285.986
R22598 a_947_1457.n0 a_947_1457.t4 282.573
R22599 a_947_1457.n1 a_947_1457.t2 202.857
R22600 a_947_1457.n1 a_947_1457.n0 173.817
R22601 a_947_1457.n1 a_947_1457.t0 20.826
R22602 a_947_1457.n2 a_947_1457.n1 20.689
R22603 a_1317_1457.t0 a_1317_1457.t1 242.857
R22604 a_1028_n2086.t0 a_1028_n2086.t1 34.8
R22605 a_4192_452.t0 a_4192_452.t1 242.857
R22606 a_2672_n271.n0 a_2672_n271.t0 358.166
R22607 a_2672_n271.t5 a_2672_n271.t3 337.399
R22608 a_2672_n271.t3 a_2672_n271.t4 285.986
R22609 a_2672_n271.n0 a_2672_n271.t5 282.573
R22610 a_2672_n271.n1 a_2672_n271.t2 202.857
R22611 a_2672_n271.n1 a_2672_n271.n0 173.817
R22612 a_2672_n271.n1 a_2672_n271.t1 20.826
R22613 a_2672_n271.n2 a_2672_n271.n1 20.689
R22614 a_2577_n286.n0 a_2577_n286.t2 362.857
R22615 a_2577_n286.t3 a_2577_n286.t4 337.399
R22616 a_2577_n286.t4 a_2577_n286.t5 298.839
R22617 a_2577_n286.n0 a_2577_n286.t3 280.405
R22618 a_2577_n286.n1 a_2577_n286.t0 200
R22619 a_2577_n286.n1 a_2577_n286.n0 172.311
R22620 a_2577_n286.n2 a_2577_n286.n1 24
R22621 a_2577_n286.n1 a_2577_n286.t1 21.212
R22622 a_6492_1216.t0 a_6492_1216.t1 242.857
R22623 a_n2677_n4116.t0 a_n2677_n4116.t1 42.707
R22624 a_7190_3666.t0 a_7190_3666.t1 242.857
R22625 a_7765_1216.t0 a_7765_1216.t1 242.857
R22626 a_4397_n30.n0 a_4397_n30.t2 358.166
R22627 a_4397_n30.t5 a_4397_n30.t4 337.399
R22628 a_4397_n30.t4 a_4397_n30.t3 285.986
R22629 a_4397_n30.n0 a_4397_n30.t5 282.573
R22630 a_4397_n30.n1 a_4397_n30.t0 202.857
R22631 a_4397_n30.n1 a_4397_n30.n0 173.817
R22632 a_4397_n30.n1 a_4397_n30.t1 20.826
R22633 a_4397_n30.n2 a_4397_n30.n1 20.689
R22634 a_4767_n30.t0 a_4767_n30.t1 242.857
R22635 a_1440_2662.t0 a_1440_2662.t1 242.857
R22636 a_865_975.t0 a_865_975.t1 242.857
R22637 ADC6_OUT[0].n0 ADC6_OUT[0].t3 1354.27
R22638 ADC6_OUT[0].n0 ADC6_OUT[0].t4 821.954
R22639 ADC6_OUT[0].n3 ADC6_OUT[0].t0 338.856
R22640 ADC6_OUT[0].n2 ADC6_OUT[0].t2 266.575
R22641 ADC6_OUT[0].n1 ADC6_OUT[0].n0 149.035
R22642 ADC6_OUT[0] ADC6_OUT[0].n3 61.785
R22643 ADC6_OUT[0].n1 ADC6_OUT[0].t1 46.723
R22644 ADC6_OUT[0].n3 ADC6_OUT[0].n2 45.176
R22645 ADC6_OUT[0].n2 ADC6_OUT[0].n1 17.317
R22646 a_6027_2928.n0 a_6027_2928.t1 362.857
R22647 a_6027_2928.t3 a_6027_2928.t4 337.399
R22648 a_6027_2928.t4 a_6027_2928.t5 298.839
R22649 a_6027_2928.n0 a_6027_2928.t3 280.405
R22650 a_6027_2928.n1 a_6027_2928.t0 200
R22651 a_6027_2928.n1 a_6027_2928.n0 172.311
R22652 a_6027_2928.n2 a_6027_2928.n1 24
R22653 a_6027_2928.n1 a_6027_2928.t2 21.212
R22654 a_4302_1924.n0 a_4302_1924.t2 362.857
R22655 a_4302_1924.t3 a_4302_1924.t5 337.399
R22656 a_4302_1924.t5 a_4302_1924.t4 298.839
R22657 a_4302_1924.n0 a_4302_1924.t3 280.405
R22658 a_4302_1924.n1 a_4302_1924.t0 200
R22659 a_4302_1924.n1 a_4302_1924.n0 172.311
R22660 a_4302_1924.n2 a_4302_1924.n1 24
R22661 a_4302_1924.n1 a_4302_1924.t1 21.212
R22662 a_5630_n5293.n0 a_5630_n5293.t0 65.063
R22663 a_5630_n5293.n0 a_5630_n5293.t2 42.011
R22664 a_5630_n5293.t1 a_5630_n5293.n0 2.113
R22665 a_9367_975.t0 a_9367_975.t1 242.857
R22666 a_3727_196.n0 a_3727_196.t0 362.857
R22667 a_3727_196.t3 a_3727_196.t5 337.399
R22668 a_3727_196.t5 a_3727_196.t4 298.839
R22669 a_3727_196.n0 a_3727_196.t3 280.405
R22670 a_3727_196.n1 a_3727_196.t1 200
R22671 a_3727_196.n1 a_3727_196.n0 172.311
R22672 a_3727_196.n2 a_3727_196.n1 24
R22673 a_3727_196.n1 a_3727_196.t2 21.212
R22674 a_3822_211.n0 a_3822_211.t2 358.166
R22675 a_3822_211.t3 a_3822_211.t5 337.399
R22676 a_3822_211.t5 a_3822_211.t4 285.986
R22677 a_3822_211.n0 a_3822_211.t3 282.573
R22678 a_3822_211.n1 a_3822_211.t0 202.857
R22679 a_3822_211.n1 a_3822_211.n0 173.817
R22680 a_3822_211.n1 a_3822_211.t1 20.826
R22681 a_3822_211.n2 a_3822_211.n1 20.689
R22682 a_2049_n6849.t0 a_2049_n6849.t1 42.707
R22683 a_2084_n6503.n0 a_2084_n6503.t0 65.064
R22684 a_2084_n6503.n0 a_2084_n6503.t2 42.011
R22685 a_2084_n6503.t1 a_2084_n6503.n0 2.113
R22686 a_3727_3651.n0 a_3727_3651.t1 362.857
R22687 a_3727_3651.t3 a_3727_3651.t4 337.399
R22688 a_3727_3651.t4 a_3727_3651.t5 298.839
R22689 a_3727_3651.n0 a_3727_3651.t3 280.405
R22690 a_3727_3651.n1 a_3727_3651.t2 200
R22691 a_3727_3651.n1 a_3727_3651.n0 172.311
R22692 a_3727_3651.n2 a_3727_3651.n1 24
R22693 a_3727_3651.n1 a_3727_3651.t0 21.212
R22694 a_2097_n30.n0 a_2097_n30.t1 358.166
R22695 a_2097_n30.t3 a_2097_n30.t5 337.399
R22696 a_2097_n30.t5 a_2097_n30.t4 285.986
R22697 a_2097_n30.n0 a_2097_n30.t3 282.573
R22698 a_2097_n30.n1 a_2097_n30.t0 202.857
R22699 a_2097_n30.n1 a_2097_n30.n0 173.817
R22700 a_2097_n30.n1 a_2097_n30.t2 20.826
R22701 a_2097_n30.n2 a_2097_n30.n1 20.689
R22702 a_2002_n45.n0 a_2002_n45.t2 362.857
R22703 a_2002_n45.t3 a_2002_n45.t5 337.399
R22704 a_2002_n45.t5 a_2002_n45.t4 298.839
R22705 a_2002_n45.n0 a_2002_n45.t3 280.405
R22706 a_2002_n45.n1 a_2002_n45.t0 200
R22707 a_2002_n45.n1 a_2002_n45.n0 172.311
R22708 a_2002_n45.n2 a_2002_n45.n1 24
R22709 a_2002_n45.n1 a_2002_n45.t1 21.212
R22710 a_5917_4445.t0 a_5917_4445.t1 242.857
R22711 a_2015_2421.t0 a_2015_2421.t1 242.857
R22712 a_3042_693.t0 a_3042_693.t1 242.857
R22713 a_2015_n271.t0 a_2015_n271.t1 242.857
R22714 a_2590_n812.t0 a_2590_n812.t1 242.857
R22715 a_6602_3651.n0 a_6602_3651.t0 362.857
R22716 a_6602_3651.t3 a_6602_3651.t5 337.399
R22717 a_6602_3651.t5 a_6602_3651.t4 298.839
R22718 a_6602_3651.n0 a_6602_3651.t3 280.405
R22719 a_6602_3651.n1 a_6602_3651.t2 200
R22720 a_6602_3651.n1 a_6602_3651.n0 172.311
R22721 a_6602_3651.n2 a_6602_3651.n1 24
R22722 a_6602_3651.n1 a_6602_3651.t1 21.212
R22723 a_5342_n1053.t0 a_5342_n1053.t1 242.857
R22724 a_3152_n286.n0 a_3152_n286.t1 362.857
R22725 a_3152_n286.t3 a_3152_n286.t4 337.399
R22726 a_3152_n286.t4 a_3152_n286.t5 298.839
R22727 a_3152_n286.n0 a_3152_n286.t3 280.405
R22728 a_3152_n286.n1 a_3152_n286.t2 200
R22729 a_3152_n286.n1 a_3152_n286.n0 172.311
R22730 a_3152_n286.n2 a_3152_n286.n1 24
R22731 a_3152_n286.n1 a_3152_n286.t0 21.212
R22732 ADC8_OUT[3].n0 ADC8_OUT[3].t4 1355.37
R22733 ADC8_OUT[3].n0 ADC8_OUT[3].t3 820.859
R22734 ADC8_OUT[3].n3 ADC8_OUT[3].t0 333.655
R22735 ADC8_OUT[3].n2 ADC8_OUT[3].t1 266.644
R22736 ADC8_OUT[3].n1 ADC8_OUT[3].n0 149.035
R22737 ADC8_OUT[3].n3 ADC8_OUT[3].n2 50.447
R22738 ADC8_OUT[3].n1 ADC8_OUT[3].t2 45.968
R22739 ADC8_OUT[3] ADC8_OUT[3].n3 22.312
R22740 ADC8_OUT[3].n2 ADC8_OUT[3].n1 17.317
R22741 a_5857_n8583.n0 a_5857_n8583.t4 1465.51
R22742 a_5857_n8583.n0 a_5857_n8583.t3 712.44
R22743 a_5857_n8583.n1 a_5857_n8583.t0 375.067
R22744 a_5857_n8583.n1 a_5857_n8583.t1 272.668
R22745 a_5857_n8583.n2 a_5857_n8583.n0 143.764
R22746 a_5857_n8583.t2 a_5857_n8583.n2 78.193
R22747 a_5857_n8583.n2 a_5857_n8583.n1 4.517
R22748 a_7067_4686.t0 a_7067_4686.t1 242.857
R22749 a_852_4671.n0 a_852_4671.t1 362.857
R22750 a_852_4671.t3 a_852_4671.t4 337.399
R22751 a_852_4671.t4 a_852_4671.t5 298.839
R22752 a_852_4671.n0 a_852_4671.t3 280.405
R22753 a_852_4671.n1 a_852_4671.t0 200
R22754 a_852_4671.n1 a_852_4671.n0 172.311
R22755 a_852_4671.n2 a_852_4671.n1 24
R22756 a_852_4671.n1 a_852_4671.t2 21.212
R22757 a_4315_4148.t0 a_4315_4148.t1 242.857
R22758 a_5465_2180.t0 a_5465_2180.t1 242.857
R22759 a_5452_437.n0 a_5452_437.t1 362.857
R22760 a_5452_437.t3 a_5452_437.t5 337.399
R22761 a_5452_437.t5 a_5452_437.t4 298.839
R22762 a_5452_437.n0 a_5452_437.t3 280.405
R22763 a_5452_437.n1 a_5452_437.t2 200
R22764 a_5452_437.n1 a_5452_437.n0 172.311
R22765 a_5452_437.n2 a_5452_437.n1 24
R22766 a_5452_437.n1 a_5452_437.t0 21.212
R22767 a_8429_n4470.t0 a_8429_n4470.t1 68.741
R22768 a_3617_3184.t0 a_3617_3184.t1 242.857
R22769 a_947_4686.n0 a_947_4686.t2 358.166
R22770 a_947_4686.t4 a_947_4686.t5 337.399
R22771 a_947_4686.t5 a_947_4686.t3 285.986
R22772 a_947_4686.n0 a_947_4686.t4 282.573
R22773 a_947_4686.n1 a_947_4686.t0 202.857
R22774 a_947_4686.n1 a_947_4686.n0 173.817
R22775 a_947_4686.n1 a_947_4686.t1 20.826
R22776 a_947_4686.n2 a_947_4686.n1 20.689
R22777 a_1317_4686.t0 a_1317_4686.t1 242.857
R22778 a_12736_n6503.n0 a_12736_n6503.t0 65.064
R22779 a_12736_n6503.n0 a_12736_n6503.t2 42.011
R22780 a_12736_n6503.t1 a_12736_n6503.n0 2.113
R22781 a_6492_4445.t0 a_6492_4445.t1 242.857
R22782 a_5342_1457.t0 a_5342_1457.t1 242.857
R22783 a_3563_n8071.n0 a_3563_n8071.t0 63.08
R22784 a_3563_n8071.n0 a_3563_n8071.t2 41.307
R22785 a_3563_n8071.t1 a_3563_n8071.n0 2.251
R22786 a_7765_4445.t0 a_7765_4445.t1 242.857
R22787 a_2049_n5092.t0 a_2049_n5092.t1 42.705
R22788 a_1522_n30.n0 a_1522_n30.t1 358.166
R22789 a_1522_n30.t4 a_1522_n30.t5 337.399
R22790 a_1522_n30.t5 a_1522_n30.t3 285.986
R22791 a_1522_n30.n0 a_1522_n30.t4 282.573
R22792 a_1522_n30.n1 a_1522_n30.t2 202.857
R22793 a_1522_n30.n1 a_1522_n30.n0 173.817
R22794 a_1522_n30.n1 a_1522_n30.t0 20.826
R22795 a_1522_n30.n2 a_1522_n30.n1 20.689
R22796 a_8902_2165.n0 a_8902_2165.t1 362.857
R22797 a_8902_2165.t5 a_8902_2165.t4 337.399
R22798 a_8902_2165.t4 a_8902_2165.t3 298.839
R22799 a_8902_2165.n0 a_8902_2165.t5 280.405
R22800 a_8902_2165.n1 a_8902_2165.t0 200
R22801 a_8902_2165.n1 a_8902_2165.n0 172.311
R22802 a_8902_2165.n2 a_8902_2165.n1 24
R22803 a_8902_2165.n1 a_8902_2165.t2 21.212
R22804 a_8915_2180.t0 a_8915_2180.t1 242.857
R22805 a_10362_n8026.n0 a_10362_n8026.t0 65.063
R22806 a_10362_n8026.n0 a_10362_n8026.t2 42.011
R22807 a_10362_n8026.t1 a_10362_n8026.n0 2.113
R22808 a_2578_n4114.t1 a_2578_n4114.t0 336.812
R22809 a_2381_n4470.n0 a_2381_n4470.t0 63.08
R22810 a_2381_n4470.n0 a_2381_n4470.t2 41.305
R22811 a_2381_n4470.t1 a_2381_n4470.n0 2.251
R22812 a_8327_1442.n0 a_8327_1442.t0 362.857
R22813 a_8327_1442.t3 a_8327_1442.t4 337.399
R22814 a_8327_1442.t4 a_8327_1442.t5 298.839
R22815 a_8327_1442.n0 a_8327_1442.t3 280.405
R22816 a_8327_1442.n1 a_8327_1442.t2 200
R22817 a_8327_1442.n1 a_8327_1442.n0 172.311
R22818 a_8327_1442.n2 a_8327_1442.n1 24
R22819 a_8327_1442.n1 a_8327_1442.t1 21.212
R22820 a_8902_678.n0 a_8902_678.t1 362.857
R22821 a_8902_678.t4 a_8902_678.t3 337.399
R22822 a_8902_678.t3 a_8902_678.t5 298.839
R22823 a_8902_678.n0 a_8902_678.t4 280.405
R22824 a_8902_678.n1 a_8902_678.t2 200
R22825 a_8902_678.n1 a_8902_678.n0 172.311
R22826 a_8902_678.n2 a_8902_678.n1 24
R22827 a_8902_678.n1 a_8902_678.t0 21.212
R22828 a_8997_693.n0 a_8997_693.t2 358.166
R22829 a_8997_693.t5 a_8997_693.t4 337.399
R22830 a_8997_693.t4 a_8997_693.t3 285.986
R22831 a_8997_693.n0 a_8997_693.t5 282.573
R22832 a_8997_693.n1 a_8997_693.t0 202.857
R22833 a_8997_693.n1 a_8997_693.n0 173.817
R22834 a_8997_693.n1 a_8997_693.t1 20.826
R22835 a_8997_693.n2 a_8997_693.n1 20.689
R22836 a_4942_n6847.t1 a_4942_n6847.t0 336.812
R22837 a_290_3184.t0 a_290_3184.t1 242.857
R22838 a_4890_n512.t0 a_4890_n512.t1 242.857
R22839 a_1892_2662.t0 a_1892_2662.t1 242.857
R22840 a_4192_3184.t0 a_4192_3184.t1 242.857
R22841 a_4767_975.t0 a_4767_975.t1 242.857
R22842 a_4972_975.n0 a_4972_975.t2 358.166
R22843 a_4972_975.t3 a_4972_975.t5 337.399
R22844 a_4972_975.t5 a_4972_975.t4 285.986
R22845 a_4972_975.n0 a_4972_975.t3 282.573
R22846 a_4972_975.n1 a_4972_975.t0 202.857
R22847 a_4972_975.n1 a_4972_975.n0 173.817
R22848 a_4972_975.n1 a_4972_975.t1 20.826
R22849 a_4972_975.n2 a_4972_975.n1 20.689
R22850 a_8422_n1053.n0 a_8422_n1053.t2 358.166
R22851 a_8422_n1053.t3 a_8422_n1053.t5 337.399
R22852 a_8422_n1053.t5 a_8422_n1053.t4 285.986
R22853 a_8422_n1053.n0 a_8422_n1053.t3 282.573
R22854 a_8422_n1053.n1 a_8422_n1053.t0 202.857
R22855 a_8422_n1053.n1 a_8422_n1053.n0 173.817
R22856 a_8422_n1053.n1 a_8422_n1053.t1 20.826
R22857 a_8422_n1053.n2 a_8422_n1053.n1 20.689
R22858 a_6040_2421.t0 a_6040_2421.t1 242.857
R22859 a_7306_n6847.t1 a_7306_n6847.t0 336.812
R22860 a_7109_n7203.n0 a_7109_n7203.t0 63.08
R22861 a_7109_n7203.n0 a_7109_n7203.t2 41.305
R22862 a_7109_n7203.t1 a_7109_n7203.n0 2.251
R22863 a_5465_3184.t0 a_5465_3184.t1 242.857
R22864 a_6040_n271.t0 a_6040_n271.t1 242.857
R22865 a_1199_n5338.n0 a_1199_n5338.t0 63.08
R22866 a_1199_n5338.n0 a_1199_n5338.t2 41.307
R22867 a_1199_n5338.t1 a_1199_n5338.n0 2.251
R22868 a_1625_n2132.n0 a_1625_n2132.t2 489.336
R22869 a_1625_n2132.n0 a_1625_n2132.t1 243.258
R22870 a_1625_n2132.t0 a_1625_n2132.n0 214.415
R22871 a_5547_n1053.n0 a_5547_n1053.t1 358.166
R22872 a_5547_n1053.t4 a_5547_n1053.t5 337.399
R22873 a_5547_n1053.t5 a_5547_n1053.t3 285.986
R22874 a_5547_n1053.n0 a_5547_n1053.t4 282.573
R22875 a_5547_n1053.n1 a_5547_n1053.t2 202.857
R22876 a_5547_n1053.n1 a_5547_n1053.n0 173.817
R22877 a_5547_n1053.n1 a_5547_n1053.t0 20.826
R22878 a_5547_n1053.n2 a_5547_n1053.n1 20.689
R22879 a_742_3907.t0 a_742_3907.t1 242.857
R22880 a_2467_2421.t0 a_2467_2421.t1 242.857
R22881 a_2467_n271.t0 a_2467_n271.t1 242.857
R22882 a_7847_n512.n0 a_7847_n512.t1 358.166
R22883 a_7847_n512.t4 a_7847_n512.t5 337.399
R22884 a_7847_n512.t5 a_7847_n512.t3 285.986
R22885 a_7847_n512.n0 a_7847_n512.t4 282.573
R22886 a_7847_n512.n1 a_7847_n512.t0 202.857
R22887 a_7847_n512.n1 a_7847_n512.n0 173.817
R22888 a_7847_n512.n1 a_7847_n512.t2 20.826
R22889 a_7847_n512.n2 a_7847_n512.n1 20.689
R22890 a_8217_n512.t0 a_8217_n512.t1 242.857
R22891 a_6697_3666.n0 a_6697_3666.t1 358.166
R22892 a_6697_3666.t3 a_6697_3666.t4 337.399
R22893 a_6697_3666.t4 a_6697_3666.t5 285.986
R22894 a_6697_3666.n0 a_6697_3666.t3 282.573
R22895 a_6697_3666.n1 a_6697_3666.t2 202.857
R22896 a_6697_3666.n1 a_6697_3666.n0 173.817
R22897 a_6697_3666.n1 a_6697_3666.t0 20.826
R22898 a_6697_3666.n2 a_6697_3666.n1 20.689
R22899 a_8340_4148.t0 a_8340_4148.t1 242.857
R22900 a_865_693.t0 a_865_693.t1 242.857
R22901 a_865_4148.t0 a_865_4148.t1 242.857
R22902 a_4890_2943.t0 a_4890_2943.t1 242.857
R22903 a_2049_n4116.t0 a_2049_n4116.t1 42.707
R22904 a_2084_n3770.n0 a_2084_n3770.t0 65.064
R22905 a_2084_n3770.n0 a_2084_n3770.t2 42.011
R22906 a_2084_n3770.t1 a_2084_n3770.n0 2.113
R22907 a_5153_n1770.t0 a_5153_n1770.t1 256.142
R22908 a_885_n1371.n1 a_885_n1371.t4 550.94
R22909 a_885_n1371.n1 a_885_n1371.t3 500.621
R22910 a_885_n1371.t2 a_885_n1371.n2 192.787
R22911 a_885_n1371.n0 a_885_n1371.t0 163.997
R22912 a_885_n1371.n2 a_885_n1371.n1 149.035
R22913 a_885_n1371.n0 a_885_n1371.t1 54.068
R22914 a_885_n1371.n2 a_885_n1371.n0 17.317
R22915 SA_OUT[1].n1 SA_OUT[1].t4 661.027
R22916 SA_OUT[1].n1 SA_OUT[1].t3 392.255
R22917 SA_OUT[1].n2 SA_OUT[1].t1 223.716
R22918 SA_OUT[1].n0 SA_OUT[1].t0 153.977
R22919 SA_OUT[1].n2 SA_OUT[1].n1 143.764
R22920 SA_OUT[1].n0 SA_OUT[1].t2 59.86
R22921 SA_OUT[1] SA_OUT[1].n3 25.019
R22922 SA_OUT[1].n3 SA_OUT[1].n0 2.258
R22923 SA_OUT[1].n3 SA_OUT[1].n2 2.258
R22924 a_4767_4148.t0 a_4767_4148.t1 242.857
R22925 a_7642_3184.t0 a_7642_3184.t1 242.857
R22926 a_8422_1457.n0 a_8422_1457.t1 358.166
R22927 a_8422_1457.t3 a_8422_1457.t5 337.399
R22928 a_8422_1457.t5 a_8422_1457.t4 285.986
R22929 a_8422_1457.n0 a_8422_1457.t3 282.573
R22930 a_8422_1457.n1 a_8422_1457.t2 202.857
R22931 a_8422_1457.n1 a_8422_1457.n0 173.817
R22932 a_8422_1457.n1 a_8422_1457.t0 20.826
R22933 a_8422_1457.n2 a_8422_1457.n1 20.689
R22934 a_9367_693.t0 a_9367_693.t1 242.857
R22935 a_5342_4686.t0 a_5342_4686.t1 242.857
R22936 a_1427_3169.n0 a_1427_3169.t1 362.857
R22937 a_1427_3169.t3 a_1427_3169.t4 337.399
R22938 a_1427_3169.t4 a_1427_3169.t5 298.839
R22939 a_1427_3169.n0 a_1427_3169.t3 280.405
R22940 a_1427_3169.n1 a_1427_3169.t0 200
R22941 a_1427_3169.n1 a_1427_3169.n0 172.311
R22942 a_1427_3169.n2 a_1427_3169.n1 24
R22943 a_1427_3169.n1 a_1427_3169.t2 21.212
R22944 a_4413_n6849.t0 a_4413_n6849.t1 42.707
R22945 a_4448_n6503.n0 a_4448_n6503.t0 65.064
R22946 a_4448_n6503.t1 a_4448_n6503.n0 42.011
R22947 a_4448_n6503.n0 a_4448_n6503.t2 2.113
R22948 a_8915_3184.t0 a_8915_3184.t1 242.857
R22949 a_3740_2180.t0 a_3740_2180.t1 242.857
R22950 a_742_n271.t0 a_742_n271.t1 242.857
R22951 a_10362_n5293.n0 a_10362_n5293.t0 65.063
R22952 a_10362_n5293.n0 a_10362_n5293.t2 42.011
R22953 a_10362_n5293.t1 a_10362_n5293.n0 2.113
R22954 a_5917_2421.t0 a_5917_2421.t1 242.857
R22955 a_n2642_n8026.n0 a_n2642_n8026.t0 65.063
R22956 a_n2642_n8026.n0 a_n2642_n8026.t2 42.011
R22957 a_n2642_n8026.t1 a_n2642_n8026.n0 2.113
R22958 a_742_3425.t0 a_742_3425.t1 242.857
R22959 a_6615_211.t0 a_6615_211.t1 242.857
R22960 a_3428_n1770.t0 a_3428_n1770.t1 256.142
R22961 a_5917_n271.t0 a_5917_n271.t1 242.857
R22962 a_902_n8026.n0 a_902_n8026.t0 65.063
R22963 a_902_n8026.n0 a_902_n8026.t2 42.011
R22964 a_902_n8026.t1 a_902_n8026.n0 2.113
R22965 a_3760_n1371.n1 a_3760_n1371.t4 550.94
R22966 a_3760_n1371.n1 a_3760_n1371.t3 500.621
R22967 a_3760_n1371.t1 a_3760_n1371.n2 192.787
R22968 a_3760_n1371.n0 a_3760_n1371.t2 163.997
R22969 a_3760_n1371.n2 a_3760_n1371.n1 149.035
R22970 a_3760_n1371.n0 a_3760_n1371.t0 54.068
R22971 a_3760_n1371.n2 a_3760_n1371.n0 17.317
R22972 SA_OUT[6].n0 SA_OUT[6].t4 661.027
R22973 SA_OUT[6].n0 SA_OUT[6].t3 392.255
R22974 SA_OUT[6].n1 SA_OUT[6].t1 223.716
R22975 SA_OUT[6].n2 SA_OUT[6].t2 153.977
R22976 SA_OUT[6].n1 SA_OUT[6].n0 143.764
R22977 SA_OUT[6].n3 SA_OUT[6].t0 58.354
R22978 SA_OUT[6] SA_OUT[6].n3 15.536
R22979 SA_OUT[6].n2 SA_OUT[6].n1 4.517
R22980 SA_OUT[6].n3 SA_OUT[6].n2 1.505
R22981 a_8327_4671.n0 a_8327_4671.t1 362.857
R22982 a_8327_4671.t3 a_8327_4671.t4 337.399
R22983 a_8327_4671.t4 a_8327_4671.t5 298.839
R22984 a_8327_4671.n0 a_8327_4671.t3 280.405
R22985 a_8327_4671.n1 a_8327_4671.t0 200
R22986 a_8327_4671.n1 a_8327_4671.n0 172.311
R22987 a_8327_4671.n2 a_8327_4671.n1 24
R22988 a_8327_4671.n1 a_8327_4671.t2 21.212
R22989 a_4315_1939.t0 a_4315_1939.t1 242.857
R22990 ADC12_OUT[3].n0 ADC12_OUT[3].t4 1355.37
R22991 ADC12_OUT[3].n0 ADC12_OUT[3].t3 820.859
R22992 ADC12_OUT[3].n3 ADC12_OUT[3].t0 322.361
R22993 ADC12_OUT[3].n2 ADC12_OUT[3].t1 266.644
R22994 ADC12_OUT[3].n1 ADC12_OUT[3].n0 149.035
R22995 ADC12_OUT[3].n3 ADC12_OUT[3].n2 61.741
R22996 ADC12_OUT[3].n1 ADC12_OUT[3].t2 45.968
R22997 ADC12_OUT[3] ADC12_OUT[3].n3 22.383
R22998 ADC12_OUT[3].n2 ADC12_OUT[3].n1 17.317
R22999 a_10589_n8583.n0 a_10589_n8583.t4 1465.51
R23000 a_10589_n8583.n0 a_10589_n8583.t3 712.44
R23001 a_10589_n8583.n1 a_10589_n8583.t0 375.067
R23002 a_10589_n8583.n1 a_10589_n8583.t1 272.668
R23003 a_10589_n8583.n2 a_10589_n8583.n0 143.764
R23004 a_10589_n8583.t2 a_10589_n8583.n2 78.193
R23005 a_10589_n8583.n2 a_10589_n8583.n1 4.517
R23006 a_6777_n4116.t0 a_6777_n4116.t1 42.707
R23007 a_7067_2662.t0 a_7067_2662.t1 242.857
R23008 a_852_2647.n0 a_852_2647.t0 362.857
R23009 a_852_2647.t3 a_852_2647.t4 337.399
R23010 a_852_2647.t4 a_852_2647.t5 298.839
R23011 a_852_2647.n0 a_852_2647.t3 280.405
R23012 a_852_2647.n1 a_852_2647.t2 200
R23013 a_852_2647.n1 a_852_2647.n0 172.311
R23014 a_852_2647.n2 a_852_2647.n1 24
R23015 a_852_2647.n1 a_852_2647.t1 21.212
R23016 a_3165_693.t0 a_3165_693.t1 242.857
R23017 a_4315_1698.t0 a_4315_1698.t1 242.857
R23018 a_12736_n3770.n0 a_12736_n3770.t0 65.064
R23019 a_12736_n3770.n0 a_12736_n3770.t2 42.011
R23020 a_12736_n3770.t1 a_12736_n3770.n0 2.113
R23021 ADC15_OUT[0].n0 ADC15_OUT[0].t3 1354.27
R23022 ADC15_OUT[0].n0 ADC15_OUT[0].t4 821.954
R23023 ADC15_OUT[0].n3 ADC15_OUT[0].t0 350.903
R23024 ADC15_OUT[0].n2 ADC15_OUT[0].t2 266.575
R23025 ADC15_OUT[0].n1 ADC15_OUT[0].n0 149.035
R23026 ADC15_OUT[0] ADC15_OUT[0].n3 61.579
R23027 ADC15_OUT[0].n1 ADC15_OUT[0].t1 46.723
R23028 ADC15_OUT[0].n3 ADC15_OUT[0].n2 33.129
R23029 ADC15_OUT[0].n2 ADC15_OUT[0].n1 17.317
R23030 a_6303_n1770.t0 a_6303_n1770.t1 256.142
R23031 SA_OUT[3].n1 SA_OUT[3].t4 661.027
R23032 SA_OUT[3].n1 SA_OUT[3].t3 392.255
R23033 SA_OUT[3].n2 SA_OUT[3].t1 223.716
R23034 SA_OUT[3].n0 SA_OUT[3].t0 153.977
R23035 SA_OUT[3].n2 SA_OUT[3].n1 143.764
R23036 SA_OUT[3].n0 SA_OUT[3].t2 59.86
R23037 SA_OUT[3] SA_OUT[3].n3 21.368
R23038 SA_OUT[3].n3 SA_OUT[3].n0 3.764
R23039 SA_OUT[3].n3 SA_OUT[3].n2 0.752
R23040 a_3042_n512.t0 a_3042_n512.t1 242.857
R23041 a_947_n812.n0 a_947_n812.t2 358.166
R23042 a_947_n812.t4 a_947_n812.t5 337.399
R23043 a_947_n812.t5 a_947_n812.t3 285.986
R23044 a_947_n812.n0 a_947_n812.t4 282.573
R23045 a_947_n812.n1 a_947_n812.t0 202.857
R23046 a_947_n812.n1 a_947_n812.n0 173.817
R23047 a_947_n812.n1 a_947_n812.t1 20.826
R23048 a_947_n812.n2 a_947_n812.n1 20.689
R23049 a_8340_452.t0 a_8340_452.t1 242.857
R23050 a_6102_n2234.n2 a_6102_n2234.t0 282.97
R23051 a_6102_n2234.n1 a_6102_n2234.t2 240.683
R23052 a_6102_n2234.n0 a_6102_n2234.t3 209.208
R23053 a_6102_n2234.n0 a_6102_n2234.t4 194.167
R23054 a_6102_n2234.t1 a_6102_n2234.n2 183.404
R23055 a_6102_n2234.n1 a_6102_n2234.n0 14.805
R23056 a_6102_n2234.n2 a_6102_n2234.n1 6.415
R23057 a_6343_n2086.t0 a_6343_n2086.t1 34.8
R23058 a_4890_693.t0 a_4890_693.t1 242.857
R23059 a_1522_3184.n0 a_1522_3184.t1 358.166
R23060 a_1522_3184.t3 a_1522_3184.t5 337.399
R23061 a_1522_3184.t5 a_1522_3184.t4 285.986
R23062 a_1522_3184.n0 a_1522_3184.t3 282.573
R23063 a_1522_3184.n1 a_1522_3184.t2 202.857
R23064 a_1522_3184.n1 a_1522_3184.n0 173.817
R23065 a_1522_3184.n1 a_1522_3184.t0 20.826
R23066 a_1522_3184.n2 a_1522_3184.n1 20.689
R23067 a_947_2662.n0 a_947_2662.t1 358.166
R23068 a_947_2662.t4 a_947_2662.t5 337.399
R23069 a_947_2662.t5 a_947_2662.t3 285.986
R23070 a_947_2662.n0 a_947_2662.t4 282.573
R23071 a_947_2662.n1 a_947_2662.t2 202.857
R23072 a_947_2662.n1 a_947_2662.n0 173.817
R23073 a_947_2662.n1 a_947_2662.t0 20.826
R23074 a_947_2662.n2 a_947_2662.n1 20.689
R23075 a_1317_2662.t0 a_1317_2662.t1 242.857
R23076 a_7752_n527.n0 a_7752_n527.t2 362.857
R23077 a_7752_n527.t3 a_7752_n527.t4 337.399
R23078 a_7752_n527.t4 a_7752_n527.t5 298.839
R23079 a_7752_n527.n0 a_7752_n527.t3 280.405
R23080 a_7752_n527.n1 a_7752_n527.t0 200
R23081 a_7752_n527.n1 a_7752_n527.n0 172.311
R23082 a_7752_n527.n2 a_7752_n527.n1 24
R23083 a_7752_n527.n1 a_7752_n527.t1 21.212
R23084 a_6492_2421.t0 a_6492_2421.t1 242.857
R23085 a_7928_n2086.t0 a_7928_n2086.t1 34.8
R23086 a_6492_n271.t0 a_6492_n271.t1 242.857
R23087 a_8488_n4114.t1 a_8488_n4114.t0 336.812
R23088 a_7765_2421.t0 a_7765_2421.t1 242.857
R23089 a_5917_211.t0 a_5917_211.t1 242.857
R23090 a_4578_n1770.n0 a_4578_n1770.t1 160.619
R23091 a_4578_n1770.t0 a_4578_n1770.n0 151.153
R23092 a_3740_1457.t0 a_3740_1457.t1 242.857
R23093 a_14131_n8026.t1 a_14131_n8026.t0 336.814
R23094 a_14072_n8071.t0 a_14072_n8071.t1 68.74
R23095 a_4942_n4114.t1 a_4942_n4114.t0 336.812
R23096 a_8422_4686.n0 a_8422_4686.t2 358.166
R23097 a_8422_4686.t3 a_8422_4686.t5 337.399
R23098 a_8422_4686.t5 a_8422_4686.t4 285.986
R23099 a_8422_4686.n0 a_8422_4686.t3 282.573
R23100 a_8422_4686.n1 a_8422_4686.t0 202.857
R23101 a_8422_4686.n1 a_8422_4686.n0 173.817
R23102 a_8422_4686.n1 a_8422_4686.t1 20.826
R23103 a_8422_4686.n2 a_8422_4686.n1 20.689
R23104 a_8792_4148.t0 a_8792_4148.t1 242.857
R23105 a_6122_211.n0 a_6122_211.t1 358.166
R23106 a_6122_211.t5 a_6122_211.t4 337.399
R23107 a_6122_211.t4 a_6122_211.t3 285.986
R23108 a_6122_211.n0 a_6122_211.t5 282.573
R23109 a_6122_211.n1 a_6122_211.t2 202.857
R23110 a_6122_211.n1 a_6122_211.n0 173.817
R23111 a_6122_211.n1 a_6122_211.t0 20.826
R23112 a_6122_211.n2 a_6122_211.n1 20.689
R23113 a_3042_2943.t0 a_3042_2943.t1 242.857
R23114 a_4767_693.t0 a_4767_693.t1 242.857
R23115 a_8915_n30.t0 a_8915_n30.t1 242.857
R23116 a_7306_n4114.t1 a_7306_n4114.t0 336.812
R23117 a_7109_n4470.n0 a_7109_n4470.t0 63.08
R23118 a_7109_n4470.n0 a_7109_n4470.t2 41.305
R23119 a_7109_n4470.t1 a_7109_n4470.n0 2.251
R23120 a_4315_1216.t0 a_4315_1216.t1 242.857
R23121 a_3810_n1770.n0 a_3810_n1770.t2 325.682
R23122 a_3810_n1770.t0 a_3810_n1770.n0 322.293
R23123 a_3810_n1770.n0 a_3810_n1770.t1 73.623
R23124 a_6492_211.t0 a_6492_211.t1 242.857
R23125 a_865_n1053.t0 a_865_n1053.t1 242.857
R23126 a_7642_452.t0 a_7642_452.t1 242.857
R23127 a_13934_n8071.n0 a_13934_n8071.t0 63.08
R23128 a_13934_n8071.n0 a_13934_n8071.t2 41.307
R23129 a_13934_n8071.t1 a_13934_n8071.n0 2.251
R23130 a_742_n812.t0 a_742_n812.t1 242.857
R23131 a_8340_1939.t0 a_8340_1939.t1 242.857
R23132 a_865_1939.t0 a_865_1939.t1 242.857
R23133 a_8792_n1053.t0 a_8792_n1053.t1 242.857
R23134 a_4397_1939.n0 a_4397_1939.t2 358.166
R23135 a_4397_1939.t4 a_4397_1939.t5 337.399
R23136 a_4397_1939.t5 a_4397_1939.t3 285.986
R23137 a_4397_1939.n0 a_4397_1939.t4 282.573
R23138 a_4397_1939.n1 a_4397_1939.t0 202.857
R23139 a_4397_1939.n1 a_4397_1939.n0 173.817
R23140 a_4397_1939.n1 a_4397_1939.t1 20.826
R23141 a_4397_1939.n2 a_4397_1939.n1 20.689
R23142 a_4767_1939.t0 a_4767_1939.t1 242.857
R23143 a_n3827_n6849.t0 a_n3827_n6849.t1 42.707
R23144 ADC13_OUT[1].n0 ADC13_OUT[1].t4 1355.37
R23145 ADC13_OUT[1].n0 ADC13_OUT[1].t3 820.859
R23146 ADC13_OUT[1].n3 ADC13_OUT[1].t0 321.608
R23147 ADC13_OUT[1].n2 ADC13_OUT[1].t1 266.644
R23148 ADC13_OUT[1].n1 ADC13_OUT[1].n0 149.035
R23149 ADC13_OUT[1].n3 ADC13_OUT[1].n2 62.494
R23150 ADC13_OUT[1] ADC13_OUT[1].n3 46.088
R23151 ADC13_OUT[1].n1 ADC13_OUT[1].t2 45.968
R23152 ADC13_OUT[1].n2 ADC13_OUT[1].n1 17.317
R23153 a_11776_n5850.n0 a_11776_n5850.t4 1465.51
R23154 a_11776_n5850.n0 a_11776_n5850.t3 712.44
R23155 a_11776_n5850.n1 a_11776_n5850.t0 375.067
R23156 a_11776_n5850.n1 a_11776_n5850.t2 272.668
R23157 a_11776_n5850.n2 a_11776_n5850.n0 143.764
R23158 a_11776_n5850.t1 a_11776_n5850.n2 78.193
R23159 a_11776_n5850.n2 a_11776_n5850.n1 4.517
R23160 a_2015_452.t0 a_2015_452.t1 242.857
R23161 a_4413_n4116.t0 a_4413_n4116.t1 42.707
R23162 a_4448_n3770.n0 a_4448_n3770.t0 65.064
R23163 a_4448_n3770.n0 a_4448_n3770.t2 42.011
R23164 a_4448_n3770.t1 a_4448_n3770.n0 2.113
R23165 a_8340_1698.t0 a_8340_1698.t1 242.857
R23166 a_865_1698.t0 a_865_1698.t1 242.857
R23167 a_n1233_n5850.n0 a_n1233_n5850.t4 1465.51
R23168 a_n1233_n5850.n0 a_n1233_n5850.t3 712.44
R23169 a_n1233_n5850.n1 a_n1233_n5850.t0 375.067
R23170 a_n1233_n5850.n1 a_n1233_n5850.t1 272.668
R23171 a_n1233_n5850.n2 a_n1233_n5850.n0 143.764
R23172 a_n1233_n5850.t2 a_n1233_n5850.n2 78.193
R23173 a_n1233_n5850.n2 a_n1233_n5850.n1 4.517
R23174 a_3740_452.t0 a_3740_452.t1 242.857
R23175 a_5342_2662.t0 a_5342_2662.t1 242.857
R23176 a_867_n4116.t0 a_867_n4116.t1 42.707
R23177 a_6122_2943.n0 a_6122_2943.t2 358.166
R23178 a_6122_2943.t3 a_6122_2943.t5 337.399
R23179 a_6122_2943.t5 a_6122_2943.t4 285.986
R23180 a_6122_2943.n0 a_6122_2943.t3 282.573
R23181 a_6122_2943.n1 a_6122_2943.t0 202.857
R23182 a_6122_2943.n1 a_6122_2943.n0 173.817
R23183 a_6122_2943.n1 a_6122_2943.t1 20.826
R23184 a_6122_2943.n2 a_6122_2943.n1 20.689
R23185 a_8327_2647.n0 a_8327_2647.t0 362.857
R23186 a_8327_2647.t3 a_8327_2647.t4 337.399
R23187 a_8327_2647.t4 a_8327_2647.t5 298.839
R23188 a_8327_2647.n0 a_8327_2647.t3 280.405
R23189 a_8327_2647.n1 a_8327_2647.t1 200
R23190 a_8327_2647.n1 a_8327_2647.n0 172.311
R23191 a_8327_2647.n2 a_8327_2647.n1 24
R23192 a_8327_2647.n1 a_8327_2647.t2 21.212
R23193 a_8792_n30.t0 a_8792_n30.t1 242.857
R23194 a_7752_4133.n0 a_7752_4133.t0 362.857
R23195 a_7752_4133.t3 a_7752_4133.t4 337.399
R23196 a_7752_4133.t4 a_7752_4133.t5 298.839
R23197 a_7752_4133.n0 a_7752_4133.t3 280.405
R23198 a_7752_4133.n1 a_7752_4133.t2 200
R23199 a_7752_4133.n1 a_7752_4133.n0 172.311
R23200 a_7752_4133.n2 a_7752_4133.n1 24
R23201 a_7752_4133.n1 a_7752_4133.t1 21.212
R23202 a_3152_960.n0 a_3152_960.t2 362.857
R23203 a_3152_960.t4 a_3152_960.t3 337.399
R23204 a_3152_960.t3 a_3152_960.t5 298.839
R23205 a_3152_960.n0 a_3152_960.t4 280.405
R23206 a_3152_960.n1 a_3152_960.t0 200
R23207 a_3152_960.n1 a_3152_960.n0 172.311
R23208 a_3152_960.n2 a_3152_960.n1 24
R23209 a_3152_960.n1 a_3152_960.t1 21.212
R23210 a_1522_211.n0 a_1522_211.t1 358.166
R23211 a_1522_211.t5 a_1522_211.t4 337.399
R23212 a_1522_211.t4 a_1522_211.t3 285.986
R23213 a_1522_211.n0 a_1522_211.t5 282.573
R23214 a_1522_211.n1 a_1522_211.t2 202.857
R23215 a_1522_211.n1 a_1522_211.n0 173.817
R23216 a_1522_211.n1 a_1522_211.t0 20.826
R23217 a_1522_211.n2 a_1522_211.n1 20.689
R23218 a_852_2928.n0 a_852_2928.t1 362.857
R23219 a_852_2928.t3 a_852_2928.t4 337.399
R23220 a_852_2928.t4 a_852_2928.t5 298.839
R23221 a_852_2928.n0 a_852_2928.t3 280.405
R23222 a_852_2928.n1 a_852_2928.t0 200
R23223 a_852_2928.n1 a_852_2928.n0 172.311
R23224 a_852_2928.n2 a_852_2928.n1 24
R23225 a_852_2928.n1 a_852_2928.t2 21.212
R23226 a_4890_3907.t0 a_4890_3907.t1 242.857
R23227 a_4972_2180.n0 a_4972_2180.t2 358.166
R23228 a_4972_2180.t3 a_4972_2180.t5 337.399
R23229 a_4972_2180.t5 a_4972_2180.t4 285.986
R23230 a_4972_2180.n0 a_4972_2180.t3 282.573
R23231 a_4972_2180.n1 a_4972_2180.t0 202.857
R23232 a_4972_2180.n1 a_4972_2180.n0 173.817
R23233 a_4972_2180.n1 a_4972_2180.t1 20.826
R23234 a_4972_2180.n2 a_4972_2180.n1 20.689
R23235 a_4877_2165.n0 a_4877_2165.t1 362.857
R23236 a_4877_2165.t4 a_4877_2165.t3 337.399
R23237 a_4877_2165.t3 a_4877_2165.t5 298.839
R23238 a_4877_2165.n0 a_4877_2165.t4 280.405
R23239 a_4877_2165.n1 a_4877_2165.t2 200
R23240 a_4877_2165.n1 a_4877_2165.n0 172.311
R23241 a_4877_2165.n2 a_4877_2165.n1 24
R23242 a_4877_2165.n1 a_4877_2165.t0 21.212
R23243 a_2590_975.t0 a_2590_975.t1 242.857
R23244 a_8997_2180.n0 a_8997_2180.t1 358.166
R23245 a_8997_2180.t4 a_8997_2180.t5 337.399
R23246 a_8997_2180.t5 a_8997_2180.t3 285.986
R23247 a_8997_2180.n0 a_8997_2180.t4 282.573
R23248 a_8997_2180.n1 a_8997_2180.t2 202.857
R23249 a_8997_2180.n1 a_8997_2180.n0 173.817
R23250 a_8997_2180.n1 a_8997_2180.t0 20.826
R23251 a_8997_2180.n2 a_8997_2180.n1 20.689
R23252 a_9367_2180.t0 a_9367_2180.t1 242.857
R23253 a_7453_n1770.n0 a_7453_n1770.t1 160.619
R23254 a_7453_n1770.t0 a_7453_n1770.n0 151.153
R23255 a_7847_4148.n0 a_7847_4148.t2 358.166
R23256 a_7847_4148.t4 a_7847_4148.t5 337.399
R23257 a_7847_4148.t5 a_7847_4148.t3 285.986
R23258 a_7847_4148.n0 a_7847_4148.t4 282.573
R23259 a_7847_4148.n1 a_7847_4148.t0 202.857
R23260 a_7847_4148.n1 a_7847_4148.n0 173.817
R23261 a_7847_4148.n1 a_7847_4148.t1 20.826
R23262 a_7847_4148.n2 a_7847_4148.n1 20.689
R23263 a_8217_4148.t0 a_8217_4148.t1 242.857
R23264 a_1892_211.t0 a_1892_211.t1 242.857
R23265 ADC9_OUT[2].n0 ADC9_OUT[2].t4 1354.27
R23266 ADC9_OUT[2].n0 ADC9_OUT[2].t3 821.954
R23267 ADC9_OUT[2].n3 ADC9_OUT[2].t0 338.103
R23268 ADC9_OUT[2].n2 ADC9_OUT[2].t1 266.575
R23269 ADC9_OUT[2].n1 ADC9_OUT[2].n0 149.035
R23270 ADC9_OUT[2].n1 ADC9_OUT[2].t2 46.723
R23271 ADC9_OUT[2].n3 ADC9_OUT[2].n2 45.929
R23272 ADC9_OUT[2] ADC9_OUT[2].n3 38.119
R23273 ADC9_OUT[2].n2 ADC9_OUT[2].n1 17.317
R23274 a_n3298_n8026.t1 a_n3298_n8026.t0 336.814
R23275 a_n3357_n8071.t0 a_n3357_n8071.t1 68.74
R23276 a_5465_3666.t0 a_5465_3666.t1 242.857
R23277 a_7190_975.t0 a_7190_975.t1 242.857
R23278 a_8792_1939.t0 a_8792_1939.t1 242.857
R23279 a_867_n7825.t0 a_867_n7825.t1 42.705
R23280 a_8422_2662.n0 a_8422_2662.t1 358.166
R23281 a_8422_2662.t3 a_8422_2662.t5 337.399
R23282 a_8422_2662.t5 a_8422_2662.t4 285.986
R23283 a_8422_2662.n0 a_8422_2662.t3 282.573
R23284 a_8422_2662.n1 a_8422_2662.t2 202.857
R23285 a_8422_2662.n1 a_8422_2662.n0 173.817
R23286 a_8422_2662.n1 a_8422_2662.t0 20.826
R23287 a_8422_2662.n2 a_8422_2662.n1 20.689
R23288 a_9178_n8026.n0 a_9178_n8026.t0 65.063
R23289 a_9178_n8026.n0 a_9178_n8026.t2 42.011
R23290 a_9178_n8026.t1 a_9178_n8026.n0 2.113
R23291 a_4890_3425.t0 a_4890_3425.t1 242.857
R23292 a_n3792_n5293.n0 a_n3792_n5293.t0 65.063
R23293 a_n3792_n5293.n0 a_n3792_n5293.t2 42.011
R23294 a_n3792_n5293.t1 a_n3792_n5293.n0 2.113
R23295 a_1427_3651.n0 a_1427_3651.t0 362.857
R23296 a_1427_3651.t3 a_1427_3651.t4 337.399
R23297 a_1427_3651.t4 a_1427_3651.t5 298.839
R23298 a_1427_3651.n0 a_1427_3651.t3 280.405
R23299 a_1427_3651.n1 a_1427_3651.t2 200
R23300 a_1427_3651.n1 a_1427_3651.n0 172.311
R23301 a_1427_3651.n2 a_1427_3651.n1 24
R23302 a_1427_3651.n1 a_1427_3651.t1 21.212
R23303 a_3617_n1053.t0 a_3617_n1053.t1 242.857
R23304 a_8603_n1770.n0 a_8603_n1770.t1 160.619
R23305 a_8603_n1770.t0 a_8603_n1770.n0 151.153
R23306 a_8915_3666.t0 a_8915_3666.t1 242.857
R23307 a_2467_n30.t0 a_2467_n30.t1 242.857
R23308 a_372_n30.n0 a_372_n30.t1 358.166
R23309 a_372_n30.t4 a_372_n30.t5 337.399
R23310 a_372_n30.t5 a_372_n30.t3 285.986
R23311 a_372_n30.n0 a_372_n30.t4 282.573
R23312 a_372_n30.n1 a_372_n30.t2 202.857
R23313 a_372_n30.n1 a_372_n30.n0 173.817
R23314 a_372_n30.n1 a_372_n30.t0 20.826
R23315 a_372_n30.n2 a_372_n30.n1 20.689
R23316 a_n1163_n8071.n0 a_n1163_n8071.t0 63.08
R23317 a_n1163_n8071.n0 a_n1163_n8071.t2 41.307
R23318 a_n1163_n8071.t1 a_n1163_n8071.n0 2.251
R23319 a_14072_n5338.t0 a_14072_n5338.t1 68.74
R23320 a_n3827_n4116.t0 a_n3827_n4116.t1 42.707
R23321 a_3152_1442.n0 a_3152_1442.t1 362.857
R23322 a_3152_1442.t3 a_3152_1442.t4 337.399
R23323 a_3152_1442.t4 a_3152_1442.t5 298.839
R23324 a_3152_1442.n0 a_3152_1442.t3 280.405
R23325 a_3152_1442.n1 a_3152_1442.t0 200
R23326 a_3152_1442.n1 a_3152_1442.n0 172.311
R23327 a_3152_1442.n2 a_3152_1442.n1 24
R23328 a_3152_1442.n1 a_3152_1442.t2 21.212
R23329 a_6040_n30.t0 a_6040_n30.t1 242.857
R23330 a_n2677_n7825.t0 a_n2677_n7825.t1 42.705
R23331 a_3042_3907.t0 a_3042_3907.t1 242.857
R23332 a_3247_1457.n0 a_3247_1457.t1 358.166
R23333 a_3247_1457.t4 a_3247_1457.t5 337.399
R23334 a_3247_1457.t5 a_3247_1457.t3 285.986
R23335 a_3247_1457.n0 a_3247_1457.t4 282.573
R23336 a_3247_1457.n1 a_3247_1457.t2 202.857
R23337 a_3247_1457.n1 a_3247_1457.n0 173.817
R23338 a_3247_1457.n1 a_3247_1457.t0 20.826
R23339 a_3247_1457.n2 a_3247_1457.n1 20.689
R23340 a_3617_1457.t0 a_3617_1457.t1 242.857
R23341 a_290_n1053.t0 a_290_n1053.t1 242.857
R23342 a_4192_n1053.t0 a_4192_n1053.t1 242.857
R23343 a_12043_n8026.t1 a_12043_n8026.t0 336.814
R23344 a_11984_n8071.t0 a_11984_n8071.t1 68.74
R23345 a_1522_3666.n0 a_1522_3666.t1 358.166
R23346 a_1522_3666.t3 a_1522_3666.t5 337.399
R23347 a_1522_3666.t5 a_1522_3666.t4 285.986
R23348 a_1522_3666.n0 a_1522_3666.t3 282.573
R23349 a_1522_3666.n1 a_1522_3666.t2 202.857
R23350 a_1522_3666.n1 a_1522_3666.n0 173.817
R23351 a_1522_3666.n1 a_1522_3666.t0 20.826
R23352 a_1522_3666.n2 a_1522_3666.n1 20.689
R23353 a_6027_3892.n0 a_6027_3892.t0 362.857
R23354 a_6027_3892.t3 a_6027_3892.t4 337.399
R23355 a_6027_3892.t4 a_6027_3892.t5 298.839
R23356 a_6027_3892.n0 a_6027_3892.t3 280.405
R23357 a_6027_3892.n1 a_6027_3892.t2 200
R23358 a_6027_3892.n1 a_6027_3892.n0 172.311
R23359 a_6027_3892.n2 a_6027_3892.n1 24
R23360 a_6027_3892.n1 a_6027_3892.t1 21.212
R23361 a_7752_196.n0 a_7752_196.t0 362.857
R23362 a_7752_196.t4 a_7752_196.t3 337.399
R23363 a_7752_196.t3 a_7752_196.t5 298.839
R23364 a_7752_196.n0 a_7752_196.t4 280.405
R23365 a_7752_196.n1 a_7752_196.t2 200
R23366 a_7752_196.n1 a_7752_196.n0 172.311
R23367 a_7752_196.n2 a_7752_196.n1 24
R23368 a_7752_196.n1 a_7752_196.t1 21.212
R23369 a_7847_211.n0 a_7847_211.t1 358.166
R23370 a_7847_211.t5 a_7847_211.t4 337.399
R23371 a_7847_211.t4 a_7847_211.t3 285.986
R23372 a_7847_211.n0 a_7847_211.t5 282.573
R23373 a_7847_211.n1 a_7847_211.t2 202.857
R23374 a_7847_211.n1 a_7847_211.n0 173.817
R23375 a_7847_211.n1 a_7847_211.t0 20.826
R23376 a_7847_211.n2 a_7847_211.n1 20.689
R23377 ADC8_OUT[1].n0 ADC8_OUT[1].t4 1355.37
R23378 ADC8_OUT[1].n0 ADC8_OUT[1].t3 820.859
R23379 ADC8_OUT[1].n3 ADC8_OUT[1].t0 328.385
R23380 ADC8_OUT[1].n2 ADC8_OUT[1].t1 266.644
R23381 ADC8_OUT[1].n1 ADC8_OUT[1].n0 149.035
R23382 ADC8_OUT[1].n3 ADC8_OUT[1].n2 55.717
R23383 ADC8_OUT[1] ADC8_OUT[1].n3 46.026
R23384 ADC8_OUT[1].n1 ADC8_OUT[1].t2 45.968
R23385 ADC8_OUT[1].n2 ADC8_OUT[1].n1 17.317
R23386 a_5857_n5850.n0 a_5857_n5850.t4 1465.51
R23387 a_5857_n5850.n0 a_5857_n5850.t3 712.44
R23388 a_5857_n5850.n1 a_5857_n5850.t0 375.067
R23389 a_5857_n5850.n1 a_5857_n5850.t2 272.668
R23390 a_5857_n5850.n2 a_5857_n5850.n0 143.764
R23391 a_5857_n5850.t1 a_5857_n5850.n2 78.193
R23392 a_5857_n5850.n2 a_5857_n5850.n1 4.517
R23393 a_6602_1924.n0 a_6602_1924.t1 362.857
R23394 a_6602_1924.t3 a_6602_1924.t5 337.399
R23395 a_6602_1924.t5 a_6602_1924.t4 298.839
R23396 a_6602_1924.n0 a_6602_1924.t3 280.405
R23397 a_6602_1924.n1 a_6602_1924.t0 200
R23398 a_6602_1924.n1 a_6602_1924.n0 172.311
R23399 a_6602_1924.n2 a_6602_1924.n1 24
R23400 a_6602_1924.n1 a_6602_1924.t2 21.212
R23401 a_8327_2928.n0 a_8327_2928.t1 362.857
R23402 a_8327_2928.t3 a_8327_2928.t4 337.399
R23403 a_8327_2928.t4 a_8327_2928.t5 298.839
R23404 a_8327_2928.n0 a_8327_2928.t3 280.405
R23405 a_8327_2928.n1 a_8327_2928.t0 200
R23406 a_8327_2928.n1 a_8327_2928.n0 172.311
R23407 a_8327_2928.n2 a_8327_2928.n1 24
R23408 a_8327_2928.n1 a_8327_2928.t2 21.212
R23409 a_1396_n8026.t1 a_1396_n8026.t0 336.814
R23410 a_1337_n8071.t0 a_1337_n8071.t1 68.74
R23411 a_5053_n2086.t0 a_5053_n2086.t1 34.8
R23412 a_290_1457.t0 a_290_1457.t1 242.857
R23413 a_7752_1683.n0 a_7752_1683.t0 362.857
R23414 a_7752_1683.t3 a_7752_1683.t4 337.399
R23415 a_7752_1683.t4 a_7752_1683.t5 298.839
R23416 a_7752_1683.n0 a_7752_1683.t3 280.405
R23417 a_7752_1683.n1 a_7752_1683.t2 200
R23418 a_7752_1683.n1 a_7752_1683.n0 172.311
R23419 a_7752_1683.n2 a_7752_1683.n1 24
R23420 a_7752_1683.n1 a_7752_1683.t1 21.212
R23421 a_4315_n271.t0 a_4315_n271.t1 242.857
R23422 ADC11_OUT[3].n0 ADC11_OUT[3].t4 1355.37
R23423 ADC11_OUT[3].n0 ADC11_OUT[3].t3 820.859
R23424 ADC11_OUT[3].n3 ADC11_OUT[3].t0 326.879
R23425 ADC11_OUT[3].n2 ADC11_OUT[3].t1 266.644
R23426 ADC11_OUT[3].n1 ADC11_OUT[3].n0 149.035
R23427 ADC11_OUT[3].n3 ADC11_OUT[3].n2 57.223
R23428 ADC11_OUT[3].n1 ADC11_OUT[3].t2 45.968
R23429 ADC11_OUT[3] ADC11_OUT[3].n3 22.446
R23430 ADC11_OUT[3].n2 ADC11_OUT[3].n1 17.317
R23431 a_4890_n812.t0 a_4890_n812.t1 242.857
R23432 a_2097_n1053.n0 a_2097_n1053.t2 358.166
R23433 a_2097_n1053.t4 a_2097_n1053.t5 337.399
R23434 a_2097_n1053.t5 a_2097_n1053.t3 285.986
R23435 a_2097_n1053.n0 a_2097_n1053.t4 282.573
R23436 a_2097_n1053.n1 a_2097_n1053.t0 202.857
R23437 a_2097_n1053.n1 a_2097_n1053.n0 173.817
R23438 a_2097_n1053.n1 a_2097_n1053.t1 20.826
R23439 a_2097_n1053.n2 a_2097_n1053.n1 20.689
R23440 a_3042_3425.t0 a_3042_3425.t1 242.857
R23441 a_4192_1457.t0 a_4192_1457.t1 242.857
R23442 a_7642_n1053.t0 a_7642_n1053.t1 242.857
R23443 a_5452_n286.n0 a_5452_n286.t1 362.857
R23444 a_5452_n286.t3 a_5452_n286.t4 337.399
R23445 a_5452_n286.t4 a_5452_n286.t5 298.839
R23446 a_5452_n286.n0 a_5452_n286.t3 280.405
R23447 a_5452_n286.n1 a_5452_n286.t2 200
R23448 a_5452_n286.n1 a_5452_n286.n0 172.311
R23449 a_5452_n286.n2 a_5452_n286.n1 24
R23450 a_5452_n286.n1 a_5452_n286.t0 21.212
R23451 a_7847_1698.n0 a_7847_1698.t2 358.166
R23452 a_7847_1698.t4 a_7847_1698.t5 337.399
R23453 a_7847_1698.t5 a_7847_1698.t3 285.986
R23454 a_7847_1698.n0 a_7847_1698.t4 282.573
R23455 a_7847_1698.n1 a_7847_1698.t0 202.857
R23456 a_7847_1698.n1 a_7847_1698.n0 173.817
R23457 a_7847_1698.n1 a_7847_1698.t1 20.826
R23458 a_7847_1698.n2 a_7847_1698.n1 20.689
R23459 a_8217_1698.t0 a_8217_1698.t1 242.857
R23460 a_7190_693.t0 a_7190_693.t1 242.857
R23461 a_3152_4671.n0 a_3152_4671.t0 362.857
R23462 a_3152_4671.t3 a_3152_4671.t4 337.399
R23463 a_3152_4671.t4 a_3152_4671.t5 298.839
R23464 a_3152_4671.n0 a_3152_4671.t3 280.405
R23465 a_3152_4671.n1 a_3152_4671.t2 200
R23466 a_3152_4671.n1 a_3152_4671.n0 172.311
R23467 a_3152_4671.n2 a_3152_4671.n1 24
R23468 a_3152_4671.n1 a_3152_4671.t1 21.212
R23469 a_6027_3410.n0 a_6027_3410.t1 362.857
R23470 a_6027_3410.t3 a_6027_3410.t4 337.399
R23471 a_6027_3410.t4 a_6027_3410.t5 298.839
R23472 a_6027_3410.n0 a_6027_3410.t3 280.405
R23473 a_6027_3410.n1 a_6027_3410.t0 200
R23474 a_6027_3410.n1 a_6027_3410.n0 172.311
R23475 a_6027_3410.n2 a_6027_3410.n1 24
R23476 a_6027_3410.n1 a_6027_3410.t2 21.212
R23477 a_7847_n812.n0 a_7847_n812.t1 358.166
R23478 a_7847_n812.t4 a_7847_n812.t5 337.399
R23479 a_7847_n812.t5 a_7847_n812.t3 285.986
R23480 a_7847_n812.n0 a_7847_n812.t4 282.573
R23481 a_7847_n812.n1 a_7847_n812.t0 202.857
R23482 a_7847_n812.n1 a_7847_n812.n0 173.817
R23483 a_7847_n812.n1 a_7847_n812.t2 20.826
R23484 a_7847_n812.n2 a_7847_n812.n1 20.689
R23485 a_8217_211.t0 a_8217_211.t1 242.857
R23486 a_3247_4686.n0 a_3247_4686.t2 358.166
R23487 a_3247_4686.t4 a_3247_4686.t5 337.399
R23488 a_3247_4686.t5 a_3247_4686.t3 285.986
R23489 a_3247_4686.n0 a_3247_4686.t4 282.573
R23490 a_3247_4686.n1 a_3247_4686.t0 202.857
R23491 a_3247_4686.n1 a_3247_4686.n0 173.817
R23492 a_3247_4686.n1 a_3247_4686.t1 20.826
R23493 a_3247_4686.n2 a_3247_4686.n1 20.689
R23494 a_3617_4686.t0 a_3617_4686.t1 242.857
R23495 a_6122_3907.n0 a_6122_3907.t1 358.166
R23496 a_6122_3907.t3 a_6122_3907.t5 337.399
R23497 a_6122_3907.t5 a_6122_3907.t4 285.986
R23498 a_6122_3907.n0 a_6122_3907.t3 282.573
R23499 a_6122_3907.n1 a_6122_3907.t2 202.857
R23500 a_6122_3907.n1 a_6122_3907.n0 173.817
R23501 a_6122_3907.n1 a_6122_3907.t0 20.826
R23502 a_6122_3907.n2 a_6122_3907.n1 20.689
R23503 a_3231_n7825.t0 a_3231_n7825.t1 42.705
R23504 a_3266_n8026.n0 a_3266_n8026.t0 65.063
R23505 a_3266_n8026.n0 a_3266_n8026.t2 42.011
R23506 a_3266_n8026.t1 a_3266_n8026.n0 2.113
R23507 a_7642_1457.t0 a_7642_1457.t1 242.857
R23508 a_7752_1201.n0 a_7752_1201.t0 362.857
R23509 a_7752_1201.t3 a_7752_1201.t4 337.399
R23510 a_7752_1201.t4 a_7752_1201.t5 298.839
R23511 a_7752_1201.n0 a_7752_1201.t3 280.405
R23512 a_7752_1201.n1 a_7752_1201.t2 200
R23513 a_7752_1201.n1 a_7752_1201.n0 172.311
R23514 a_7752_1201.n2 a_7752_1201.n1 24
R23515 a_7752_1201.n1 a_7752_1201.t1 21.212
R23516 a_2753_n2086.t0 a_2753_n2086.t1 34.8
R23517 a_3231_n6849.t0 a_3231_n6849.t1 42.707
R23518 a_7847_1216.n0 a_7847_1216.t2 358.166
R23519 a_7847_1216.t4 a_7847_1216.t5 337.399
R23520 a_7847_1216.t5 a_7847_1216.t3 285.986
R23521 a_7847_1216.n0 a_7847_1216.t4 282.573
R23522 a_7847_1216.n1 a_7847_1216.t0 202.857
R23523 a_7847_1216.n1 a_7847_1216.n0 173.817
R23524 a_7847_1216.n1 a_7847_1216.t1 20.826
R23525 a_7847_1216.n2 a_7847_1216.n1 20.689
R23526 a_8217_1216.t0 a_8217_1216.t1 242.857
R23527 a_7177_n45.n0 a_7177_n45.t2 362.857
R23528 a_7177_n45.t4 a_7177_n45.t3 337.399
R23529 a_7177_n45.t3 a_7177_n45.t5 298.839
R23530 a_7177_n45.n0 a_7177_n45.t4 280.405
R23531 a_7177_n45.n1 a_7177_n45.t0 200
R23532 a_7177_n45.n1 a_7177_n45.n0 172.311
R23533 a_7177_n45.n2 a_7177_n45.n1 24
R23534 a_7177_n45.n1 a_7177_n45.t1 21.212
R23535 a_n314_n4378.n3 a_n314_n4378.t3 475.39
R23536 a_n314_n4378.n3 a_n314_n4378.n2 255.792
R23537 a_n314_n4378.t4 a_n314_n4378.t6 228.696
R23538 a_n314_n4378.n2 a_n314_n4378.t2 185.704
R23539 a_n314_n4378.n0 a_n314_n4378.t4 126.761
R23540 a_n314_n4378.n1 a_n314_n4378.t5 126.284
R23541 a_n314_n4378.n1 a_n314_n4378.t1 126.284
R23542 a_n314_n4378.t0 a_n314_n4378.n3 124.375
R23543 a_n314_n4378.t1 a_n314_n4378.n0 115.122
R23544 a_n314_n4378.n0 a_n314_n4378.t7 111.229
R23545 a_n314_n4378.n2 a_n314_n4378.n1 8.764
R23546 a_290_4686.t0 a_290_4686.t1 242.857
R23547 a_1317_n512.t0 a_1317_n512.t1 242.857
R23548 a_4192_4686.t0 a_4192_4686.t1 242.857
R23549 a_6122_3425.n0 a_6122_3425.t2 358.166
R23550 a_6122_3425.t3 a_6122_3425.t5 337.399
R23551 a_6122_3425.t5 a_6122_3425.t4 285.986
R23552 a_6122_3425.n0 a_6122_3425.t3 282.573
R23553 a_6122_3425.n1 a_6122_3425.t0 202.857
R23554 a_6122_3425.n1 a_6122_3425.n0 173.817
R23555 a_6122_3425.n1 a_6122_3425.t1 20.826
R23556 a_6122_3425.n2 a_6122_3425.n1 20.689
R23557 a_1440_4148.t0 a_1440_4148.t1 242.857
R23558 a_7765_3184.t0 a_7765_3184.t1 242.857
R23559 a_2590_2180.t0 a_2590_2180.t1 242.857
R23560 a_8340_n271.t0 a_8340_n271.t1 242.857
R23561 a_742_975.t0 a_742_975.t1 242.857
R23562 a_865_n271.t0 a_865_n271.t1 242.857
R23563 a_3042_n812.t0 a_3042_n812.t1 242.857
R23564 a_n2345_n7203.n0 a_n2345_n7203.t0 63.08
R23565 a_n2345_n7203.n0 a_n2345_n7203.t2 41.305
R23566 a_n2345_n7203.t1 a_n2345_n7203.n0 2.251
R23567 a_3903_n2086.t0 a_3903_n2086.t1 34.8
R23568 a_4877_437.n0 a_4877_437.t2 362.857
R23569 a_4877_437.t4 a_4877_437.t3 337.399
R23570 a_4877_437.t3 a_4877_437.t5 298.839
R23571 a_4877_437.n0 a_4877_437.t4 280.405
R23572 a_4877_437.n1 a_4877_437.t0 200
R23573 a_4877_437.n1 a_4877_437.n0 172.311
R23574 a_4877_437.n2 a_4877_437.n1 24
R23575 a_4877_437.n1 a_4877_437.t1 21.212
R23576 a_4972_452.n0 a_4972_452.t1 358.166
R23577 a_4972_452.t5 a_4972_452.t4 337.399
R23578 a_4972_452.t4 a_4972_452.t3 285.986
R23579 a_4972_452.n0 a_4972_452.t5 282.573
R23580 a_4972_452.n1 a_4972_452.t2 202.857
R23581 a_4972_452.n1 a_4972_452.n0 173.817
R23582 a_4972_452.n1 a_4972_452.t0 20.826
R23583 a_4972_452.n2 a_4972_452.n1 20.689
R23584 a_4767_n271.t0 a_4767_n271.t1 242.857
R23585 a_2590_693.t0 a_2590_693.t1 242.857
R23586 a_7752_n827.n0 a_7752_n827.t2 362.857
R23587 a_7752_n827.t3 a_7752_n827.t4 337.399
R23588 a_7752_n827.t4 a_7752_n827.t5 298.839
R23589 a_7752_n827.n0 a_7752_n827.t3 280.405
R23590 a_7752_n827.n1 a_7752_n827.t0 200
R23591 a_7752_n827.n1 a_7752_n827.n0 172.311
R23592 a_7752_n827.n2 a_7752_n827.n1 24
R23593 a_7752_n827.n1 a_7752_n827.t1 21.212
R23594 a_3165_1939.t0 a_3165_1939.t1 242.857
R23595 a_947_2943.n0 a_947_2943.t2 358.166
R23596 a_947_2943.t4 a_947_2943.t5 337.399
R23597 a_947_2943.t5 a_947_2943.t3 285.986
R23598 a_947_2943.n0 a_947_2943.t4 282.573
R23599 a_947_2943.n1 a_947_2943.t0 202.857
R23600 a_947_2943.n1 a_947_2943.n0 173.817
R23601 a_947_2943.n1 a_947_2943.t1 20.826
R23602 a_947_2943.n2 a_947_2943.n1 20.689
R23603 a_1317_2943.t0 a_1317_2943.t1 242.857
R23604 a_7642_4686.t0 a_7642_4686.t1 242.857
R23605 a_3617_211.t0 a_3617_211.t1 242.857
R23606 ADC12_OUT[1].n0 ADC12_OUT[1].t4 1355.37
R23607 ADC12_OUT[1].n0 ADC12_OUT[1].t3 820.859
R23608 ADC12_OUT[1].n3 ADC12_OUT[1].t0 328.385
R23609 ADC12_OUT[1].n2 ADC12_OUT[1].t1 266.644
R23610 ADC12_OUT[1].n1 ADC12_OUT[1].n0 149.035
R23611 ADC12_OUT[1].n3 ADC12_OUT[1].n2 55.717
R23612 ADC12_OUT[1] ADC12_OUT[1].n3 45.972
R23613 ADC12_OUT[1].n1 ADC12_OUT[1].t2 45.968
R23614 ADC12_OUT[1].n2 ADC12_OUT[1].n1 17.317
R23615 a_10589_n5850.n0 a_10589_n5850.t4 1465.51
R23616 a_10589_n5850.n0 a_10589_n5850.t3 712.44
R23617 a_10589_n5850.n1 a_10589_n5850.t0 375.067
R23618 a_10589_n5850.n1 a_10589_n5850.t2 272.668
R23619 a_10589_n5850.n2 a_10589_n5850.n0 143.764
R23620 a_10589_n5850.t1 a_10589_n5850.n2 78.193
R23621 a_10589_n5850.n2 a_10589_n5850.n1 4.517
R23622 a_935_n1770.n0 a_935_n1770.t2 322.294
R23623 a_935_n1770.n1 a_935_n1770.n0 229.466
R23624 a_935_n1770.t0 a_935_n1770.n1 151.15
R23625 a_935_n1770.n0 a_935_n1770.t1 73.623
R23626 a_3760_n8026.t1 a_3760_n8026.t0 336.814
R23627 a_3701_n8071.t0 a_3701_n8071.t1 68.74
R23628 a_7752_4430.n0 a_7752_4430.t0 362.857
R23629 a_7752_4430.t3 a_7752_4430.t4 337.399
R23630 a_7752_4430.t4 a_7752_4430.t5 298.839
R23631 a_7752_4430.n0 a_7752_4430.t3 280.405
R23632 a_7752_4430.n1 a_7752_4430.t2 200
R23633 a_7752_4430.n1 a_7752_4430.n0 172.311
R23634 a_7752_4430.n2 a_7752_4430.n1 24
R23635 a_7752_4430.n1 a_7752_4430.t1 21.212
R23636 a_1892_n1053.t0 a_1892_n1053.t1 242.857
R23637 ADC1_OUT[0].n0 ADC1_OUT[0].t3 1354.27
R23638 ADC1_OUT[0].n0 ADC1_OUT[0].t4 821.954
R23639 ADC1_OUT[0].n3 ADC1_OUT[0].t0 351.656
R23640 ADC1_OUT[0].n2 ADC1_OUT[0].t2 266.575
R23641 ADC1_OUT[0].n1 ADC1_OUT[0].n0 149.035
R23642 ADC1_OUT[0] ADC1_OUT[0].n3 61.651
R23643 ADC1_OUT[0].n1 ADC1_OUT[0].t1 46.723
R23644 ADC1_OUT[0].n3 ADC1_OUT[0].n2 32.376
R23645 ADC1_OUT[0].n2 ADC1_OUT[0].n1 17.317
R23646 a_6124_n8026.t1 a_6124_n8026.t0 336.814
R23647 a_6065_n8071.t0 a_6065_n8071.t1 68.74
R23648 a_852_n45.n0 a_852_n45.t2 362.857
R23649 a_852_n45.t4 a_852_n45.t3 337.399
R23650 a_852_n45.t3 a_852_n45.t5 298.839
R23651 a_852_n45.n0 a_852_n45.t4 280.405
R23652 a_852_n45.n1 a_852_n45.t0 200
R23653 a_852_n45.n1 a_852_n45.n0 172.311
R23654 a_852_n45.n2 a_852_n45.n1 24
R23655 a_852_n45.n1 a_852_n45.t1 21.212
R23656 a_7847_4445.n0 a_7847_4445.t1 358.166
R23657 a_7847_4445.t4 a_7847_4445.t5 337.399
R23658 a_7847_4445.t5 a_7847_4445.t3 285.986
R23659 a_7847_4445.n0 a_7847_4445.t4 282.573
R23660 a_7847_4445.n1 a_7847_4445.t2 202.857
R23661 a_7847_4445.n1 a_7847_4445.n0 173.817
R23662 a_7847_4445.n1 a_7847_4445.t0 20.826
R23663 a_7847_4445.n2 a_7847_4445.n1 20.689
R23664 a_8217_4445.t0 a_8217_4445.t1 242.857
R23665 a_6615_1939.t0 a_6615_1939.t1 242.857
R23666 a_5342_452.t0 a_5342_452.t1 242.857
R23667 a_6110_n1770.n0 a_6110_n1770.t2 325.682
R23668 a_6110_n1770.t0 a_6110_n1770.n0 322.293
R23669 a_6110_n1770.n0 a_6110_n1770.t1 73.623
R23670 a_6152_n1770.t0 a_6152_n1770.t1 213.924
R23671 a_3152_2647.n0 a_3152_2647.t1 362.857
R23672 a_3152_2647.t3 a_3152_2647.t4 337.399
R23673 a_3152_2647.t4 a_3152_2647.t5 298.839
R23674 a_3152_2647.n0 a_3152_2647.t3 280.405
R23675 a_3152_2647.n1 a_3152_2647.t2 200
R23676 a_3152_2647.n1 a_3152_2647.n0 172.311
R23677 a_3152_2647.n2 a_3152_2647.n1 24
R23678 a_3152_2647.n1 a_3152_2647.t0 21.212
R23679 a_5342_n512.t0 a_5342_n512.t1 242.857
R23680 a_1337_n5338.t0 a_1337_n5338.t1 68.74
R23681 a_n3827_n5092.t0 a_n3827_n5092.t1 42.705
R23682 a_3247_2662.n0 a_3247_2662.t2 358.166
R23683 a_3247_2662.t4 a_3247_2662.t5 337.399
R23684 a_3247_2662.t5 a_3247_2662.t3 285.986
R23685 a_3247_2662.n0 a_3247_2662.t4 282.573
R23686 a_3247_2662.n1 a_3247_2662.t0 202.857
R23687 a_3247_2662.n1 a_3247_2662.n0 173.817
R23688 a_3247_2662.n1 a_3247_2662.t1 20.826
R23689 a_3247_2662.n2 a_3247_2662.n1 20.689
R23690 a_3617_2662.t0 a_3617_2662.t1 242.857
R23691 a_4413_n5092.t0 a_4413_n5092.t1 42.705
R23692 a_11846_n5338.n0 a_11846_n5338.t0 63.08
R23693 a_11846_n5338.n0 a_11846_n5338.t2 41.307
R23694 a_11846_n5338.t1 a_11846_n5338.n0 2.251
R23695 a_1892_4148.t0 a_1892_4148.t1 242.857
R23696 a_8792_n271.t0 a_8792_n271.t1 242.857
R23697 ADC6_OUT[2].n0 ADC6_OUT[2].t4 1354.27
R23698 ADC6_OUT[2].n0 ADC6_OUT[2].t3 821.954
R23699 ADC6_OUT[2].n3 ADC6_OUT[2].t0 341.115
R23700 ADC6_OUT[2].n2 ADC6_OUT[2].t1 266.575
R23701 ADC6_OUT[2].n1 ADC6_OUT[2].n0 149.035
R23702 ADC6_OUT[2].n1 ADC6_OUT[2].t2 46.723
R23703 ADC6_OUT[2].n3 ADC6_OUT[2].n2 42.917
R23704 ADC6_OUT[2] ADC6_OUT[2].n3 38.066
R23705 ADC6_OUT[2].n2 ADC6_OUT[2].n1 17.317
R23706 a_3493_n7216.n0 a_3493_n7216.t4 1464.36
R23707 a_3493_n7216.n0 a_3493_n7216.t3 713.588
R23708 a_3493_n7216.n1 a_3493_n7216.t2 374.998
R23709 a_3493_n7216.n1 a_3493_n7216.t1 273.351
R23710 a_3493_n7216.n2 a_3493_n7216.n0 143.764
R23711 a_3493_n7216.t0 a_3493_n7216.n2 78.209
R23712 a_3493_n7216.n2 a_3493_n7216.n1 4.517
R23713 a_9027_n1770.t0 a_9027_n1770.t1 213.924
R23714 a_5917_n30.t0 a_5917_n30.t1 242.857
R23715 a_7190_1939.t0 a_7190_1939.t1 242.857
R23716 a_n1460_n5293.n0 a_n1460_n5293.t0 65.063
R23717 a_n1460_n5293.n0 a_n1460_n5293.t2 42.011
R23718 a_n1460_n5293.t1 a_n1460_n5293.n0 2.113
R23719 ADC5_OUT[0].n0 ADC5_OUT[0].t3 1354.27
R23720 ADC5_OUT[0].n0 ADC5_OUT[0].t4 821.954
R23721 ADC5_OUT[0].n3 ADC5_OUT[0].t0 349.397
R23722 ADC5_OUT[0].n2 ADC5_OUT[0].t1 266.575
R23723 ADC5_OUT[0].n1 ADC5_OUT[0].n0 149.035
R23724 ADC5_OUT[0] ADC5_OUT[0].n3 61.561
R23725 ADC5_OUT[0].n1 ADC5_OUT[0].t2 46.723
R23726 ADC5_OUT[0].n3 ADC5_OUT[0].n2 34.635
R23727 ADC5_OUT[0].n2 ADC5_OUT[0].n1 17.317
R23728 a_290_975.t0 a_290_975.t1 242.857
R23729 a_2610_n1371.n1 a_2610_n1371.t4 550.94
R23730 a_2610_n1371.n1 a_2610_n1371.t3 500.621
R23731 a_2610_n1371.t2 a_2610_n1371.n2 192.787
R23732 a_2610_n1371.n0 a_2610_n1371.t0 163.997
R23733 a_2610_n1371.n2 a_2610_n1371.n1 149.035
R23734 a_2610_n1371.n0 a_2610_n1371.t1 54.068
R23735 a_2610_n1371.n2 a_2610_n1371.n0 17.317
R23736 SA_OUT[4].n1 SA_OUT[4].t4 661.027
R23737 SA_OUT[4].n1 SA_OUT[4].t3 392.255
R23738 SA_OUT[4].n2 SA_OUT[4].t1 223.716
R23739 SA_OUT[4].n0 SA_OUT[4].t2 153.977
R23740 SA_OUT[4].n2 SA_OUT[4].n1 143.764
R23741 SA_OUT[4].n0 SA_OUT[4].t0 59.86
R23742 SA_OUT[4] SA_OUT[4].n3 19.535
R23743 SA_OUT[4].n3 SA_OUT[4].n0 2.258
R23744 SA_OUT[4].n3 SA_OUT[4].n2 2.258
R23745 a_5342_2943.t0 a_5342_2943.t1 242.857
R23746 a_290_2662.t0 a_290_2662.t1 242.857
R23747 a_13602_n7825.t0 a_13602_n7825.t1 42.705
R23748 a_13637_n8026.n0 a_13637_n8026.t0 65.063
R23749 a_13637_n8026.n0 a_13637_n8026.t2 42.011
R23750 a_13637_n8026.t1 a_13637_n8026.n0 2.113
R23751 a_4192_2662.t0 a_4192_2662.t1 242.857
R23752 a_4315_975.t0 a_4315_975.t1 242.857
R23753 ADC3_OUT[3].n0 ADC3_OUT[3].t4 1355.37
R23754 ADC3_OUT[3].n0 ADC3_OUT[3].t3 820.859
R23755 ADC3_OUT[3].n3 ADC3_OUT[3].t0 326.879
R23756 ADC3_OUT[3].n2 ADC3_OUT[3].t2 266.644
R23757 ADC3_OUT[3].n1 ADC3_OUT[3].n0 149.035
R23758 ADC3_OUT[3].n3 ADC3_OUT[3].n2 57.223
R23759 ADC3_OUT[3].n1 ADC3_OUT[3].t1 45.968
R23760 ADC3_OUT[3] ADC3_OUT[3].n3 22.08
R23761 ADC3_OUT[3].n2 ADC3_OUT[3].n1 17.317
R23762 a_n2345_n4470.n0 a_n2345_n4470.t0 63.08
R23763 a_n2345_n4470.n0 a_n2345_n4470.t2 41.305
R23764 a_n2345_n4470.t1 a_n2345_n4470.n0 2.251
R23765 a_1440_1698.t0 a_1440_1698.t1 242.857
R23766 a_8993_n2422.n3 a_8993_n2422.t3 475.39
R23767 a_8993_n2422.t4 a_8993_n2422.t6 228.696
R23768 a_8993_n2422.n2 a_8993_n2422.t2 185.704
R23769 a_8993_n2422.n3 a_8993_n2422.n2 165.472
R23770 a_8993_n2422.n0 a_8993_n2422.t4 126.761
R23771 a_8993_n2422.n1 a_8993_n2422.t5 126.284
R23772 a_8993_n2422.n1 a_8993_n2422.t1 126.284
R23773 a_8993_n2422.t0 a_8993_n2422.n3 124.375
R23774 a_8993_n2422.t1 a_8993_n2422.n0 115.122
R23775 a_8993_n2422.n0 a_8993_n2422.t7 111.229
R23776 a_8993_n2422.n2 a_8993_n2422.n1 8.764
R23777 a_13602_n6849.t0 a_13602_n6849.t1 42.707
R23778 a_2015_1457.t0 a_2015_1457.t1 242.857
R23779 a_7642_2662.t0 a_7642_2662.t1 242.857
R23780 a_2578_n5293.t1 a_2578_n5293.t0 336.814
R23781 a_7067_4148.t0 a_7067_4148.t1 242.857
R23782 a_7752_2406.n0 a_7752_2406.t0 362.857
R23783 a_7752_2406.t3 a_7752_2406.t4 337.399
R23784 a_7752_2406.t4 a_7752_2406.t5 298.839
R23785 a_7752_2406.n0 a_7752_2406.t3 280.405
R23786 a_7752_2406.n1 a_7752_2406.t2 200
R23787 a_7752_2406.n1 a_7752_2406.n0 172.311
R23788 a_7752_2406.n2 a_7752_2406.n1 24
R23789 a_7752_2406.n1 a_7752_2406.t1 21.212
R23790 a_n2415_n7216.n0 a_n2415_n7216.t4 1464.36
R23791 a_n2415_n7216.n0 a_n2415_n7216.t3 713.588
R23792 a_n2415_n7216.n1 a_n2415_n7216.t0 374.998
R23793 a_n2415_n7216.n1 a_n2415_n7216.t1 273.351
R23794 a_n2415_n7216.n2 a_n2415_n7216.n0 143.764
R23795 a_n2415_n7216.t2 a_n2415_n7216.n2 78.209
R23796 a_n2415_n7216.n2 a_n2415_n7216.n1 4.517
R23797 a_1440_1216.t0 a_1440_1216.t1 242.857
R23798 a_8422_2943.n0 a_8422_2943.t2 358.166
R23799 a_8422_2943.t3 a_8422_2943.t5 337.399
R23800 a_8422_2943.t5 a_8422_2943.t4 285.986
R23801 a_8422_2943.n0 a_8422_2943.t3 282.573
R23802 a_8422_2943.n1 a_8422_2943.t0 202.857
R23803 a_8422_2943.n1 a_8422_2943.n0 173.817
R23804 a_8422_2943.n1 a_8422_2943.t1 20.826
R23805 a_8422_2943.n2 a_8422_2943.n1 20.689
R23806 a_7847_2421.n0 a_7847_2421.t2 358.166
R23807 a_7847_2421.t4 a_7847_2421.t5 337.399
R23808 a_7847_2421.t5 a_7847_2421.t3 285.986
R23809 a_7847_2421.n0 a_7847_2421.t4 282.573
R23810 a_7847_2421.n1 a_7847_2421.t0 202.857
R23811 a_7847_2421.n1 a_7847_2421.n0 173.817
R23812 a_7847_2421.n1 a_7847_2421.t1 20.826
R23813 a_7847_2421.n2 a_7847_2421.n1 20.689
R23814 a_8217_2421.t0 a_8217_2421.t1 242.857
R23815 a_1129_n7216.n0 a_1129_n7216.t4 1464.36
R23816 a_1129_n7216.n0 a_1129_n7216.t3 713.588
R23817 a_1129_n7216.n1 a_1129_n7216.t0 374.998
R23818 a_1129_n7216.n1 a_1129_n7216.t1 273.351
R23819 a_1129_n7216.n2 a_1129_n7216.n0 143.764
R23820 a_1129_n7216.t2 a_1129_n7216.n2 78.209
R23821 a_1129_n7216.n2 a_1129_n7216.n1 4.517
R23822 a_852_3892.n0 a_852_3892.t0 362.857
R23823 a_852_3892.t3 a_852_3892.t4 337.399
R23824 a_852_3892.t4 a_852_3892.t5 298.839
R23825 a_852_3892.n0 a_852_3892.t3 280.405
R23826 a_852_3892.n1 a_852_3892.t2 200
R23827 a_852_3892.n1 a_852_3892.n0 172.311
R23828 a_852_3892.n2 a_852_3892.n1 24
R23829 a_852_3892.n1 a_852_3892.t1 21.212
R23830 a_3152_2928.n0 a_3152_2928.t1 362.857
R23831 a_3152_2928.t3 a_3152_2928.t4 337.399
R23832 a_3152_2928.t4 a_3152_2928.t5 298.839
R23833 a_3152_2928.n0 a_3152_2928.t3 280.405
R23834 a_3152_2928.n1 a_3152_2928.t0 200
R23835 a_3152_2928.n1 a_3152_2928.n0 172.311
R23836 a_3152_2928.n2 a_3152_2928.n1 24
R23837 a_3152_2928.n1 a_3152_2928.t2 21.212
R23838 a_12736_n5293.n0 a_12736_n5293.t0 65.063
R23839 a_12736_n5293.n0 a_12736_n5293.t2 42.011
R23840 a_12736_n5293.t1 a_12736_n5293.n0 2.113
R23841 a_4890_975.t0 a_4890_975.t1 242.857
R23842 a_6040_n1053.t0 a_6040_n1053.t1 242.857
R23843 a_3701_n5338.t0 a_3701_n5338.t1 68.74
R23844 a_947_3907.n0 a_947_3907.t2 358.166
R23845 a_947_3907.t4 a_947_3907.t5 337.399
R23846 a_947_3907.t5 a_947_3907.t3 285.986
R23847 a_947_3907.n0 a_947_3907.t4 282.573
R23848 a_947_3907.n1 a_947_3907.t0 202.857
R23849 a_947_3907.n1 a_947_3907.n0 173.817
R23850 a_947_3907.n1 a_947_3907.t1 20.826
R23851 a_947_3907.n2 a_947_3907.n1 20.689
R23852 a_1317_3907.t0 a_1317_3907.t1 242.857
R23853 a_4192_975.t0 a_4192_975.t1 242.857
R23854 a_902_n6503.n0 a_902_n6503.t0 65.064
R23855 a_902_n6503.t1 a_902_n6503.n0 42.011
R23856 a_902_n6503.n0 a_902_n6503.t2 2.113
R23857 a_742_2180.t0 a_742_2180.t1 242.857
R23858 a_2467_n1053.t0 a_2467_n1053.t1 242.857
R23859 a_5927_n5338.n0 a_5927_n5338.t0 63.08
R23860 a_5927_n5338.n0 a_5927_n5338.t2 41.307
R23861 a_5927_n5338.t1 a_5927_n5338.n0 2.251
R23862 a_6065_n5338.t0 a_6065_n5338.t1 68.74
R23863 a_7765_3666.t0 a_7765_3666.t1 242.857
R23864 a_6697_1939.n0 a_6697_1939.t2 358.166
R23865 a_6697_1939.t3 a_6697_1939.t4 337.399
R23866 a_6697_1939.t4 a_6697_1939.t5 285.986
R23867 a_6697_1939.n0 a_6697_1939.t3 282.573
R23868 a_6697_1939.n1 a_6697_1939.t0 202.857
R23869 a_6697_1939.n1 a_6697_1939.n0 173.817
R23870 a_6697_1939.n1 a_6697_1939.t1 20.826
R23871 a_6697_1939.n2 a_6697_1939.n1 20.689
R23872 a_2015_4686.t0 a_2015_4686.t1 242.857
R23873 a_1892_1698.t0 a_1892_1698.t1 242.857
R23874 a_1427_1924.n0 a_1427_1924.t0 362.857
R23875 a_1427_1924.t3 a_1427_1924.t4 337.399
R23876 a_1427_1924.t4 a_1427_1924.t5 298.839
R23877 a_1427_1924.n0 a_1427_1924.t3 280.405
R23878 a_1427_1924.n1 a_1427_1924.t2 200
R23879 a_1427_1924.n1 a_1427_1924.n0 172.311
R23880 a_1427_1924.n2 a_1427_1924.n1 24
R23881 a_1427_1924.n1 a_1427_1924.t1 21.212
R23882 a_2002_1442.n0 a_2002_1442.t1 362.857
R23883 a_2002_1442.t3 a_2002_1442.t5 337.399
R23884 a_2002_1442.t5 a_2002_1442.t4 298.839
R23885 a_2002_1442.n0 a_2002_1442.t3 280.405
R23886 a_2002_1442.n1 a_2002_1442.t0 200
R23887 a_2002_1442.n1 a_2002_1442.n0 172.311
R23888 a_2002_1442.n2 a_2002_1442.n1 24
R23889 a_2002_1442.n1 a_2002_1442.t2 21.212
R23890 a_852_3410.n0 a_852_3410.t1 362.857
R23891 a_852_3410.t3 a_852_3410.t4 337.399
R23892 a_852_3410.t4 a_852_3410.t5 298.839
R23893 a_852_3410.n0 a_852_3410.t3 280.405
R23894 a_852_3410.n1 a_852_3410.t0 200
R23895 a_852_3410.n1 a_852_3410.n0 172.311
R23896 a_852_3410.n2 a_852_3410.n1 24
R23897 a_852_3410.n1 a_852_3410.t2 21.212
R23898 a_290_693.t0 a_290_693.t1 242.857
R23899 a_6040_1457.t0 a_6040_1457.t1 242.857
R23900 a_947_3425.n0 a_947_3425.t2 358.166
R23901 a_947_3425.t4 a_947_3425.t5 337.399
R23902 a_947_3425.t5 a_947_3425.t3 285.986
R23903 a_947_3425.n0 a_947_3425.t4 282.573
R23904 a_947_3425.n1 a_947_3425.t0 202.857
R23905 a_947_3425.n1 a_947_3425.n0 173.817
R23906 a_947_3425.n1 a_947_3425.t1 20.826
R23907 a_947_3425.n2 a_947_3425.n1 20.689
R23908 a_1317_3425.t0 a_1317_3425.t1 242.857
R23909 a_2097_1457.n0 a_2097_1457.t1 358.166
R23910 a_2097_1457.t4 a_2097_1457.t5 337.399
R23911 a_2097_1457.t5 a_2097_1457.t3 285.986
R23912 a_2097_1457.n0 a_2097_1457.t4 282.573
R23913 a_2097_1457.n1 a_2097_1457.t2 202.857
R23914 a_2097_1457.n1 a_2097_1457.n0 173.817
R23915 a_2097_1457.n1 a_2097_1457.t0 20.826
R23916 a_2097_1457.n2 a_2097_1457.n1 20.689
R23917 a_2467_1457.t0 a_2467_1457.t1 242.857
R23918 a_5917_n1053.t0 a_5917_n1053.t1 242.857
R23919 a_4315_693.t0 a_4315_693.t1 242.857
R23920 a_1440_4445.t0 a_1440_4445.t1 242.857
R23921 a_3727_n286.n0 a_3727_n286.t2 362.857
R23922 a_3727_n286.t3 a_3727_n286.t4 337.399
R23923 a_3727_n286.t4 a_3727_n286.t5 298.839
R23924 a_3727_n286.n0 a_3727_n286.t3 280.405
R23925 a_3727_n286.n1 a_3727_n286.t0 200
R23926 a_3727_n286.n1 a_3727_n286.n0 172.311
R23927 a_3727_n286.n2 a_3727_n286.n1 24
R23928 a_3727_n286.n1 a_3727_n286.t1 21.212
R23929 a_3822_n271.n0 a_3822_n271.t2 358.166
R23930 a_3822_n271.t5 a_3822_n271.t4 337.399
R23931 a_3822_n271.t4 a_3822_n271.t3 285.986
R23932 a_3822_n271.n0 a_3822_n271.t5 282.573
R23933 a_3822_n271.n1 a_3822_n271.t0 202.857
R23934 a_3822_n271.n1 a_3822_n271.n0 173.817
R23935 a_3822_n271.n1 a_3822_n271.t1 20.826
R23936 a_3822_n271.n2 a_3822_n271.n1 20.689
R23937 a_6040_211.t0 a_6040_211.t1 242.857
R23938 ADC15_OUT[2].n0 ADC15_OUT[2].t4 1354.27
R23939 ADC15_OUT[2].n0 ADC15_OUT[2].t3 821.954
R23940 ADC15_OUT[2].n3 ADC15_OUT[2].t0 337.35
R23941 ADC15_OUT[2].n2 ADC15_OUT[2].t1 266.575
R23942 ADC15_OUT[2].n1 ADC15_OUT[2].n0 149.035
R23943 ADC15_OUT[2].n1 ADC15_OUT[2].t2 46.723
R23944 ADC15_OUT[2].n3 ADC15_OUT[2].n2 46.682
R23945 ADC15_OUT[2] ADC15_OUT[2].n3 38.065
R23946 ADC15_OUT[2].n2 ADC15_OUT[2].n1 17.317
R23947 a_13864_n7216.n0 a_13864_n7216.t4 1464.36
R23948 a_13864_n7216.n0 a_13864_n7216.t3 713.588
R23949 a_13864_n7216.n1 a_13864_n7216.t0 374.998
R23950 a_13864_n7216.n1 a_13864_n7216.t2 273.351
R23951 a_13864_n7216.n2 a_13864_n7216.n0 143.764
R23952 a_13864_n7216.t1 a_13864_n7216.n2 78.209
R23953 a_13864_n7216.n2 a_13864_n7216.n1 4.517
R23954 a_13033_n8071.n0 a_13033_n8071.t0 63.08
R23955 a_13033_n8071.n0 a_13033_n8071.t2 41.307
R23956 a_13033_n8071.t1 a_13033_n8071.n0 2.251
R23957 a_5452_1442.n0 a_5452_1442.t2 362.857
R23958 a_5452_1442.t3 a_5452_1442.t4 337.399
R23959 a_5452_1442.t4 a_5452_1442.t5 298.839
R23960 a_5452_1442.n0 a_5452_1442.t3 280.405
R23961 a_5452_1442.n1 a_5452_1442.t0 200
R23962 a_5452_1442.n1 a_5452_1442.n0 172.311
R23963 a_5452_1442.n2 a_5452_1442.n1 24
R23964 a_5452_1442.n1 a_5452_1442.t1 21.212
R23965 a_1892_1216.t0 a_1892_1216.t1 242.857
R23966 a_7765_n30.t0 a_7765_n30.t1 242.857
R23967 a_5342_3907.t0 a_5342_3907.t1 242.857
R23968 a_5547_1457.n0 a_5547_1457.t1 358.166
R23969 a_5547_1457.t4 a_5547_1457.t5 337.399
R23970 a_5547_1457.t5 a_5547_1457.t3 285.986
R23971 a_5547_1457.n0 a_5547_1457.t4 282.573
R23972 a_5547_1457.n1 a_5547_1457.t2 202.857
R23973 a_5547_1457.n1 a_5547_1457.n0 173.817
R23974 a_5547_1457.n1 a_5547_1457.t0 20.826
R23975 a_5547_1457.n2 a_5547_1457.n1 20.689
R23976 a_5917_1457.t0 a_5917_1457.t1 242.857
R23977 a_3165_n271.t0 a_3165_n271.t1 242.857
R23978 a_2311_n5850.n0 a_2311_n5850.t4 1465.51
R23979 a_2311_n5850.n0 a_2311_n5850.t3 712.44
R23980 a_2311_n5850.n1 a_2311_n5850.t0 375.067
R23981 a_2311_n5850.n1 a_2311_n5850.t1 272.668
R23982 a_2311_n5850.n2 a_2311_n5850.n0 143.764
R23983 a_2311_n5850.t2 a_2311_n5850.n2 78.193
R23984 a_2311_n5850.n2 a_2311_n5850.n1 4.517
R23985 a_4942_n5293.t1 a_4942_n5293.t0 336.814
R23986 a_6492_n1053.t0 a_6492_n1053.t1 242.857
R23987 ADC11_OUT[1].n0 ADC11_OUT[1].t4 1355.37
R23988 ADC11_OUT[1].n0 ADC11_OUT[1].t3 820.859
R23989 ADC11_OUT[1].n3 ADC11_OUT[1].t0 333.655
R23990 ADC11_OUT[1].n2 ADC11_OUT[1].t2 266.644
R23991 ADC11_OUT[1].n1 ADC11_OUT[1].n0 149.035
R23992 ADC11_OUT[1].n3 ADC11_OUT[1].n2 50.447
R23993 ADC11_OUT[1] ADC11_OUT[1].n3 46.026
R23994 ADC11_OUT[1].n1 ADC11_OUT[1].t1 45.968
R23995 ADC11_OUT[1].n2 ADC11_OUT[1].n1 17.317
R23996 a_2002_4671.n0 a_2002_4671.t0 362.857
R23997 a_2002_4671.t3 a_2002_4671.t5 337.399
R23998 a_2002_4671.t5 a_2002_4671.t4 298.839
R23999 a_2002_4671.n0 a_2002_4671.t3 280.405
R24000 a_2002_4671.n1 a_2002_4671.t2 200
R24001 a_2002_4671.n1 a_2002_4671.n0 172.311
R24002 a_2002_4671.n2 a_2002_4671.n1 24
R24003 a_2002_4671.n1 a_2002_4671.t1 21.212
R24004 a_7067_1698.t0 a_7067_1698.t1 242.857
R24005 a_7306_n5293.t1 a_7306_n5293.t0 336.814
R24006 a_8327_3892.n0 a_8327_3892.t0 362.857
R24007 a_8327_3892.t3 a_8327_3892.t4 337.399
R24008 a_8327_3892.t4 a_8327_3892.t5 298.839
R24009 a_8327_3892.n0 a_8327_3892.t3 280.405
R24010 a_8327_3892.n1 a_8327_3892.t2 200
R24011 a_8327_3892.n1 a_8327_3892.n0 172.311
R24012 a_8327_3892.n2 a_8327_3892.n1 24
R24013 a_8327_3892.n1 a_8327_3892.t1 21.212
R24014 a_6040_4686.t0 a_6040_4686.t1 242.857
R24015 a_11846_n8071.n0 a_11846_n8071.t0 63.08
R24016 a_11846_n8071.n0 a_11846_n8071.t2 41.307
R24017 a_11846_n8071.t1 a_11846_n8071.n0 2.251
R24018 a_2097_4686.n0 a_2097_4686.t1 358.166
R24019 a_2097_4686.t4 a_2097_4686.t5 337.399
R24020 a_2097_4686.t5 a_2097_4686.t3 285.986
R24021 a_2097_4686.n0 a_2097_4686.t4 282.573
R24022 a_2097_4686.n1 a_2097_4686.t2 202.857
R24023 a_2097_4686.n1 a_2097_4686.n0 173.817
R24024 a_2097_4686.n1 a_2097_4686.t0 20.826
R24025 a_2097_4686.n2 a_2097_4686.n1 20.689
R24026 a_2467_4686.t0 a_2467_4686.t1 242.857
R24027 a_11514_n7825.t0 a_11514_n7825.t1 42.705
R24028 a_902_n3770.n0 a_902_n3770.t0 65.064
R24029 a_902_n3770.n0 a_902_n3770.t2 42.011
R24030 a_902_n3770.t1 a_902_n3770.n0 2.113
R24031 a_4192_693.t0 a_4192_693.t1 242.857
R24032 a_8340_n30.t0 a_8340_n30.t1 242.857
R24033 a_6615_n271.t0 a_6615_n271.t1 242.857
R24034 a_5342_3425.t0 a_5342_3425.t1 242.857
R24035 a_6492_1457.t0 a_6492_1457.t1 242.857
R24036 a_1317_n812.t0 a_1317_n812.t1 242.857
R24037 a_1199_n8071.n0 a_1199_n8071.t0 63.08
R24038 a_1199_n8071.n0 a_1199_n8071.t2 41.307
R24039 a_1199_n8071.t1 a_1199_n8071.n0 2.251
R24040 a_11514_n6849.t1 a_11514_n6849.t0 42.707
R24041 a_215_n8026.t1 a_215_n8026.t0 336.814
R24042 a_156_n8071.t0 a_156_n8071.t1 68.74
R24043 a_5452_4671.n0 a_5452_4671.t0 362.857
R24044 a_5452_4671.t3 a_5452_4671.t4 337.399
R24045 a_5452_4671.t4 a_5452_4671.t5 298.839
R24046 a_5452_4671.n0 a_5452_4671.t3 280.405
R24047 a_5452_4671.n1 a_5452_4671.t2 200
R24048 a_5452_4671.n1 a_5452_4671.n0 172.311
R24049 a_5452_4671.n2 a_5452_4671.n1 24
R24050 a_5452_4671.n1 a_5452_4671.t1 21.212
R24051 a_8902_4133.n0 a_8902_4133.t1 362.857
R24052 a_8902_4133.t5 a_8902_4133.t4 337.399
R24053 a_8902_4133.t4 a_8902_4133.t3 298.839
R24054 a_8902_4133.n0 a_8902_4133.t5 280.405
R24055 a_8902_4133.n1 a_8902_4133.t0 200
R24056 a_8902_4133.n1 a_8902_4133.n0 172.311
R24057 a_8902_4133.n2 a_8902_4133.n1 24
R24058 a_8902_4133.n1 a_8902_4133.t2 21.212
R24059 a_1440_211.t0 a_1440_211.t1 242.857
R24060 a_1892_4445.t0 a_1892_4445.t1 242.857
R24061 a_7067_1216.t0 a_7067_1216.t1 242.857
R24062 a_8327_3410.n0 a_8327_3410.t1 362.857
R24063 a_8327_3410.t3 a_8327_3410.t4 337.399
R24064 a_8327_3410.t4 a_8327_3410.t5 298.839
R24065 a_8327_3410.n0 a_8327_3410.t3 280.405
R24066 a_8327_3410.n1 a_8327_3410.t0 200
R24067 a_8327_3410.n1 a_8327_3410.n0 172.311
R24068 a_8327_3410.n2 a_8327_3410.n1 24
R24069 a_8327_3410.n1 a_8327_3410.t2 21.212
R24070 a_9143_n7825.t0 a_9143_n7825.t1 42.705
R24071 a_7039_n4483.n0 a_7039_n4483.t3 1464.36
R24072 a_7039_n4483.n0 a_7039_n4483.t4 713.588
R24073 a_7039_n4483.n1 a_7039_n4483.t0 374.998
R24074 a_7039_n4483.n1 a_7039_n4483.t2 273.351
R24075 a_7039_n4483.n2 a_7039_n4483.n0 143.764
R24076 a_7039_n4483.t1 a_7039_n4483.n2 78.209
R24077 a_7039_n4483.n2 a_7039_n4483.n1 4.517
R24078 a_8217_n30.t0 a_8217_n30.t1 242.857
R24079 a_5547_4686.n0 a_5547_4686.t1 358.166
R24080 a_5547_4686.t4 a_5547_4686.t5 337.399
R24081 a_5547_4686.t5 a_5547_4686.t3 285.986
R24082 a_5547_4686.n0 a_5547_4686.t4 282.573
R24083 a_5547_4686.n1 a_5547_4686.t2 202.857
R24084 a_5547_4686.n1 a_5547_4686.n0 173.817
R24085 a_5547_4686.n1 a_5547_4686.t0 20.826
R24086 a_5547_4686.n2 a_5547_4686.n1 20.689
R24087 a_5917_4686.t0 a_5917_4686.t1 242.857
R24088 a_8422_3907.n0 a_8422_3907.t1 358.166
R24089 a_8422_3907.t3 a_8422_3907.t5 337.399
R24090 a_8422_3907.t5 a_8422_3907.t4 285.986
R24091 a_8422_3907.n0 a_8422_3907.t3 282.573
R24092 a_8422_3907.n1 a_8422_3907.t2 202.857
R24093 a_8422_3907.n1 a_8422_3907.n0 173.817
R24094 a_8422_3907.n1 a_8422_3907.t0 20.826
R24095 a_8422_3907.n2 a_8422_3907.n1 20.689
R24096 a_3740_n30.t0 a_3740_n30.t1 242.857
R24097 a_2015_2662.t0 a_2015_2662.t1 242.857
R24098 a_6602_196.n0 a_6602_196.t0 362.857
R24099 a_6602_196.t3 a_6602_196.t5 337.399
R24100 a_6602_196.t5 a_6602_196.t4 298.839
R24101 a_6602_196.n0 a_6602_196.t3 280.405
R24102 a_6602_196.n1 a_6602_196.t1 200
R24103 a_6602_196.n1 a_6602_196.n0 172.311
R24104 a_6602_196.n2 a_6602_196.n1 24
R24105 a_6602_196.n1 a_6602_196.t2 21.212
R24106 a_6697_211.n0 a_6697_211.t2 358.166
R24107 a_6697_211.t4 a_6697_211.t3 337.399
R24108 a_6697_211.t3 a_6697_211.t5 285.986
R24109 a_6697_211.n0 a_6697_211.t4 282.573
R24110 a_6697_211.n1 a_6697_211.t0 202.857
R24111 a_6697_211.n1 a_6697_211.n0 173.817
R24112 a_6697_211.n1 a_6697_211.t1 20.826
R24113 a_6697_211.n2 a_6697_211.n1 20.689
R24114 a_7190_n271.t0 a_7190_n271.t1 242.857
R24115 a_10659_n5338.n0 a_10659_n5338.t0 63.08
R24116 a_10659_n5338.n0 a_10659_n5338.t2 41.307
R24117 a_10659_n5338.t1 a_10659_n5338.n0 2.251
R24118 a_8997_n512.n0 a_8997_n512.t2 358.166
R24119 a_8997_n512.t4 a_8997_n512.t5 337.399
R24120 a_8997_n512.t5 a_8997_n512.t3 285.986
R24121 a_8997_n512.n0 a_8997_n512.t4 282.573
R24122 a_8997_n512.n1 a_8997_n512.t0 202.857
R24123 a_8997_n512.n1 a_8997_n512.n0 173.817
R24124 a_8997_n512.n1 a_8997_n512.t1 20.826
R24125 a_8997_n512.n2 a_8997_n512.n1 20.689
R24126 a_1440_2421.t0 a_1440_2421.t1 242.857
R24127 a_2519_n7203.t0 a_2519_n7203.t1 68.741
R24128 a_2015_n30.t0 a_2015_n30.t1 242.857
R24129 a_2127_n1770.t0 a_2127_n1770.n0 182.779
R24130 a_2127_n1770.n0 a_2127_n1770.t1 111.474
R24131 Din[10].n0 Din[10].t0 215.292
R24132 Din[10].n0 Din[10].t1 187.376
R24133 Din[10] Din[10].n0 84.894
R24134 a_3617_n512.t0 a_3617_n512.t1 242.857
R24135 a_6492_4686.t0 a_6492_4686.t1 242.857
R24136 a_8422_3425.n0 a_8422_3425.t1 358.166
R24137 a_8422_3425.t3 a_8422_3425.t5 337.399
R24138 a_8422_3425.t5 a_8422_3425.t4 285.986
R24139 a_8422_3425.n0 a_8422_3425.t3 282.573
R24140 a_8422_3425.n1 a_8422_3425.t2 202.857
R24141 a_8422_3425.n1 a_8422_3425.n0 173.817
R24142 a_8422_3425.n1 a_8422_3425.t0 20.826
R24143 a_8422_3425.n2 a_8422_3425.n1 20.689
R24144 a_4890_2180.t0 a_4890_2180.t1 242.857
R24145 a_3740_4148.t0 a_3740_4148.t1 242.857
R24146 a_6778_n2086.t0 a_6778_n2086.t1 34.8
R24147 ADC10_OUT[3].n0 ADC10_OUT[3].t4 1355.37
R24148 ADC10_OUT[3].n0 ADC10_OUT[3].t3 820.859
R24149 ADC10_OUT[3].n3 ADC10_OUT[3].t0 327.632
R24150 ADC10_OUT[3].n2 ADC10_OUT[3].t2 266.644
R24151 ADC10_OUT[3].n1 ADC10_OUT[3].n0 149.035
R24152 ADC10_OUT[3].n3 ADC10_OUT[3].n2 56.47
R24153 ADC10_OUT[3].n1 ADC10_OUT[3].t1 45.968
R24154 ADC10_OUT[3] ADC10_OUT[3].n3 22.382
R24155 ADC10_OUT[3].n2 ADC10_OUT[3].n1 17.317
R24156 a_5342_n812.t0 a_5342_n812.t1 242.857
R24157 a_7067_4445.t0 a_7067_4445.t1 242.857
R24158 a_n966_n6847.t1 a_n966_n6847.t0 336.812
R24159 a_5465_1939.t0 a_5465_1939.t1 242.857
R24160 a_n2642_n6503.n0 a_n2642_n6503.t0 65.064
R24161 a_n2642_n6503.n0 a_n2642_n6503.t2 42.011
R24162 a_n2642_n6503.t1 a_n2642_n6503.n0 2.113
R24163 a_3247_2943.n0 a_3247_2943.t2 358.166
R24164 a_3247_2943.t4 a_3247_2943.t5 337.399
R24165 a_3247_2943.t5 a_3247_2943.t3 285.986
R24166 a_3247_2943.n0 a_3247_2943.t4 282.573
R24167 a_3247_2943.n1 a_3247_2943.t0 202.857
R24168 a_3247_2943.n1 a_3247_2943.n0 173.817
R24169 a_3247_2943.n1 a_3247_2943.t1 20.826
R24170 a_3247_2943.n2 a_3247_2943.n1 20.689
R24171 a_3617_2943.t0 a_3617_2943.t1 242.857
R24172 a_2002_2647.n0 a_2002_2647.t0 362.857
R24173 a_2002_2647.t3 a_2002_2647.t5 337.399
R24174 a_2002_2647.t5 a_2002_2647.t4 298.839
R24175 a_2002_2647.n0 a_2002_2647.t3 280.405
R24176 a_2002_2647.n1 a_2002_2647.t2 200
R24177 a_2002_2647.n1 a_2002_2647.n0 172.311
R24178 a_2002_2647.n2 a_2002_2647.n1 24
R24179 a_2002_2647.n1 a_2002_2647.t1 21.212
R24180 a_290_n512.t0 a_290_n512.t1 242.857
R24181 a_6040_2662.t0 a_6040_2662.t1 242.857
R24182 a_4192_n512.t0 a_4192_n512.t1 242.857
R24183 Din[12].n0 Din[12].t0 215.292
R24184 Din[12].n0 Din[12].t1 187.376
R24185 Din[12] Din[12].n0 84.912
R24186 a_7252_n2234.n2 a_7252_n2234.t1 282.97
R24187 a_7252_n2234.n1 a_7252_n2234.t4 240.683
R24188 a_7252_n2234.n0 a_7252_n2234.t2 209.208
R24189 a_7252_n2234.n0 a_7252_n2234.t3 194.167
R24190 a_7252_n2234.t0 a_7252_n2234.n2 183.404
R24191 a_7252_n2234.n1 a_7252_n2234.n0 14.805
R24192 a_7252_n2234.n2 a_7252_n2234.n1 6.415
R24193 a_7642_975.t0 a_7642_975.t1 242.857
R24194 a_2097_2662.n0 a_2097_2662.t1 358.166
R24195 a_2097_2662.t4 a_2097_2662.t5 337.399
R24196 a_2097_2662.t5 a_2097_2662.t3 285.986
R24197 a_2097_2662.n0 a_2097_2662.t4 282.573
R24198 a_2097_2662.n1 a_2097_2662.t2 202.857
R24199 a_2097_2662.n1 a_2097_2662.n0 173.817
R24200 a_2097_2662.n1 a_2097_2662.t0 20.826
R24201 a_2097_2662.n2 a_2097_2662.n1 20.689
R24202 a_2467_2662.t0 a_2467_2662.t1 242.857
R24203 a_8902_n527.n0 a_8902_n527.t2 362.857
R24204 a_8902_n527.t5 a_8902_n527.t4 337.399
R24205 a_8902_n527.t4 a_8902_n527.t3 298.839
R24206 a_8902_n527.n0 a_8902_n527.t5 280.405
R24207 a_8902_n527.n1 a_8902_n527.t0 200
R24208 a_8902_n527.n1 a_8902_n527.n0 172.311
R24209 a_8902_n527.n2 a_8902_n527.n1 24
R24210 a_8902_n527.n1 a_8902_n527.t1 21.212
R24211 a_7765_211.t0 a_7765_211.t1 242.857
R24212 a_8915_1939.t0 a_8915_1939.t1 242.857
R24213 a_2002_437.n0 a_2002_437.t1 362.857
R24214 a_2002_437.t3 a_2002_437.t5 337.399
R24215 a_2002_437.t5 a_2002_437.t4 298.839
R24216 a_2002_437.n0 a_2002_437.t3 280.405
R24217 a_2002_437.n1 a_2002_437.t2 200
R24218 a_2002_437.n1 a_2002_437.n0 172.311
R24219 a_2002_437.n2 a_2002_437.n1 24
R24220 a_2002_437.n1 a_2002_437.t0 21.212
R24221 a_5927_n8071.n0 a_5927_n8071.t0 63.08
R24222 a_5927_n8071.n0 a_5927_n8071.t2 41.307
R24223 a_5927_n8071.t1 a_5927_n8071.n0 2.251
R24224 a_290_2943.t0 a_290_2943.t1 242.857
R24225 a_7752_3169.n0 a_7752_3169.t0 362.857
R24226 a_7752_3169.t3 a_7752_3169.t4 337.399
R24227 a_7752_3169.t4 a_7752_3169.t5 298.839
R24228 a_7752_3169.n0 a_7752_3169.t3 280.405
R24229 a_7752_3169.n1 a_7752_3169.t2 200
R24230 a_7752_3169.n1 a_7752_3169.n0 172.311
R24231 a_7752_3169.n2 a_7752_3169.n1 24
R24232 a_7752_3169.n1 a_7752_3169.t1 21.212
R24233 a_1892_2421.t0 a_1892_2421.t1 242.857
R24234 a_8902_1683.n0 a_8902_1683.t1 362.857
R24235 a_8902_1683.t5 a_8902_1683.t4 337.399
R24236 a_8902_1683.t4 a_8902_1683.t3 298.839
R24237 a_8902_1683.n0 a_8902_1683.t5 280.405
R24238 a_8902_1683.n1 a_8902_1683.t0 200
R24239 a_8902_1683.n1 a_8902_1683.n0 172.311
R24240 a_8902_1683.n2 a_8902_1683.n1 24
R24241 a_8902_1683.n1 a_8902_1683.t2 21.212
R24242 a_4192_2943.t0 a_4192_2943.t1 242.857
R24243 a_5595_n7825.t0 a_5595_n7825.t1 42.705
R24244 a_7642_n512.t0 a_7642_n512.t1 242.857
R24245 a_5547_2662.n0 a_5547_2662.t1 358.166
R24246 a_5547_2662.t4 a_5547_2662.t5 337.399
R24247 a_5547_2662.t5 a_5547_2662.t3 285.986
R24248 a_5547_2662.n0 a_5547_2662.t4 282.573
R24249 a_5547_2662.n1 a_5547_2662.t2 202.857
R24250 a_5547_2662.n1 a_5547_2662.n0 173.817
R24251 a_5547_2662.n1 a_5547_2662.t0 20.826
R24252 a_5547_2662.n2 a_5547_2662.n1 20.689
R24253 a_5917_2662.t0 a_5917_2662.t1 242.857
R24254 a_7847_3184.n0 a_7847_3184.t2 358.166
R24255 a_7847_3184.t4 a_7847_3184.t5 337.399
R24256 a_7847_3184.t5 a_7847_3184.t3 285.986
R24257 a_7847_3184.n0 a_7847_3184.t4 282.573
R24258 a_7847_3184.n1 a_7847_3184.t0 202.857
R24259 a_7847_3184.n1 a_7847_3184.n0 173.817
R24260 a_7847_3184.n1 a_7847_3184.t1 20.826
R24261 a_7847_3184.n2 a_7847_3184.n1 20.689
R24262 a_8217_3184.t0 a_8217_3184.t1 242.857
R24263 a_3042_2180.t0 a_3042_2180.t1 242.857
R24264 a_5595_n6849.t1 a_5595_n6849.t0 42.707
R24265 a_7190_n1053.t0 a_7190_n1053.t1 242.857
R24266 a_5002_n1770.t0 a_5002_n1770.t1 213.924
R24267 a_n1163_n5338.n0 a_n1163_n5338.t0 63.08
R24268 a_n1163_n5338.n0 a_n1163_n5338.t2 41.307
R24269 a_n1163_n5338.t1 a_n1163_n5338.n0 2.251
R24270 a_n1025_n5338.t0 a_n1025_n5338.t1 68.74
R24271 ADC9_OUT[0].n0 ADC9_OUT[0].t3 1354.27
R24272 ADC9_OUT[0].n0 ADC9_OUT[0].t4 821.954
R24273 ADC9_OUT[0].n3 ADC9_OUT[0].t0 346.385
R24274 ADC9_OUT[0].n2 ADC9_OUT[0].t2 266.575
R24275 ADC9_OUT[0].n1 ADC9_OUT[0].n0 149.035
R24276 ADC9_OUT[0] ADC9_OUT[0].n3 61.704
R24277 ADC9_OUT[0].n1 ADC9_OUT[0].t1 46.723
R24278 ADC9_OUT[0].n3 ADC9_OUT[0].n2 37.647
R24279 ADC9_OUT[0].n2 ADC9_OUT[0].n1 17.317
R24280 a_18_n5338.n0 a_18_n5338.t0 63.08
R24281 a_18_n5338.n0 a_18_n5338.t2 41.307
R24282 a_18_n5338.t1 a_18_n5338.n0 2.251
R24283 a_156_n5338.t0 a_156_n5338.t1 68.74
R24284 ADC3_OUT[1].n0 ADC3_OUT[1].t4 1355.37
R24285 ADC3_OUT[1].n0 ADC3_OUT[1].t3 820.859
R24286 ADC3_OUT[1].n3 ADC3_OUT[1].t0 329.138
R24287 ADC3_OUT[1].n2 ADC3_OUT[1].t1 266.644
R24288 ADC3_OUT[1].n1 ADC3_OUT[1].n0 149.035
R24289 ADC3_OUT[1].n3 ADC3_OUT[1].n2 54.964
R24290 ADC3_OUT[1].n1 ADC3_OUT[1].t2 45.968
R24291 ADC3_OUT[1] ADC3_OUT[1].n3 45.74
R24292 ADC3_OUT[1].n2 ADC3_OUT[1].n1 17.317
R24293 a_1522_1939.n0 a_1522_1939.t1 358.166
R24294 a_1522_1939.t3 a_1522_1939.t5 337.399
R24295 a_1522_1939.t5 a_1522_1939.t4 285.986
R24296 a_1522_1939.n0 a_1522_1939.t3 282.573
R24297 a_1522_1939.n1 a_1522_1939.t2 202.857
R24298 a_1522_1939.n1 a_1522_1939.n0 173.817
R24299 a_1522_1939.n1 a_1522_1939.t0 20.826
R24300 a_1522_1939.n2 a_1522_1939.n1 20.689
R24301 a_4883_n7203.t0 a_4883_n7203.t1 68.741
R24302 a_7642_2943.t0 a_7642_2943.t1 242.857
R24303 a_1317_975.t0 a_1317_975.t1 242.857
R24304 a_5465_n1053.t0 a_5465_n1053.t1 242.857
R24305 a_8902_1201.n0 a_8902_1201.t1 362.857
R24306 a_8902_1201.t5 a_8902_1201.t4 337.399
R24307 a_8902_1201.t4 a_8902_1201.t3 298.839
R24308 a_8902_1201.n0 a_8902_1201.t5 280.405
R24309 a_8902_1201.n1 a_8902_1201.t0 200
R24310 a_8902_1201.n1 a_8902_1201.n0 172.311
R24311 a_8902_1201.n2 a_8902_1201.n1 24
R24312 a_8902_1201.n1 a_8902_1201.t2 21.212
R24313 a_4315_n1053.t0 a_4315_n1053.t1 242.857
R24314 a_7247_n7203.t0 a_7247_n7203.t1 68.741
R24315 a_4960_n1770.n0 a_4960_n1770.t1 322.294
R24316 a_4960_n1770.n1 a_4960_n1770.n0 229.466
R24317 a_4960_n1770.t0 a_4960_n1770.n1 151.15
R24318 a_4960_n1770.n0 a_4960_n1770.t2 73.623
R24319 a_6492_2662.t0 a_6492_2662.t1 242.857
R24320 a_n966_n4114.t1 a_n966_n4114.t0 336.812
R24321 a_3740_1698.t0 a_3740_1698.t1 242.857
R24322 a_n2642_n3770.n0 a_n2642_n3770.t0 65.064
R24323 a_n2642_n3770.n0 a_n2642_n3770.t2 42.011
R24324 a_n2642_n3770.t1 a_n2642_n3770.n0 2.113
R24325 a_8340_n1053.t0 a_8340_n1053.t1 242.857
R24326 a_7067_2421.t0 a_7067_2421.t1 242.857
R24327 a_3165_452.t0 a_3165_452.t1 242.857
R24328 a_9672_n8026.t1 a_9672_n8026.t0 336.814
R24329 a_9613_n8071.t0 a_9613_n8071.t1 68.74
R24330 a_7877_n1770.t0 a_7877_n1770.t1 213.924
R24331 a_4315_1457.t0 a_4315_1457.t1 242.857
R24332 a_2002_2928.n0 a_2002_2928.t1 362.857
R24333 a_2002_2928.t3 a_2002_2928.t5 337.399
R24334 a_2002_2928.t5 a_2002_2928.t4 298.839
R24335 a_2002_2928.n0 a_2002_2928.t3 280.405
R24336 a_2002_2928.n1 a_2002_2928.t0 200
R24337 a_2002_2928.n1 a_2002_2928.n0 172.311
R24338 a_2002_2928.n2 a_2002_2928.n1 24
R24339 a_2002_2928.n1 a_2002_2928.t2 21.212
R24340 a_6122_2180.n0 a_6122_2180.t2 358.166
R24341 a_6122_2180.t3 a_6122_2180.t5 337.399
R24342 a_6122_2180.t5 a_6122_2180.t4 285.986
R24343 a_6122_2180.n0 a_6122_2180.t3 282.573
R24344 a_6122_2180.n1 a_6122_2180.t0 202.857
R24345 a_6122_2180.n1 a_6122_2180.n0 173.817
R24346 a_6122_2180.n1 a_6122_2180.t1 20.826
R24347 a_6122_2180.n2 a_6122_2180.n1 20.689
R24348 a_4972_4148.n0 a_4972_4148.t2 358.166
R24349 a_4972_4148.t3 a_4972_4148.t5 337.399
R24350 a_4972_4148.t5 a_4972_4148.t4 285.986
R24351 a_4972_4148.n0 a_4972_4148.t3 282.573
R24352 a_4972_4148.n1 a_4972_4148.t0 202.857
R24353 a_4972_4148.n1 a_4972_4148.n0 173.817
R24354 a_4972_4148.n1 a_4972_4148.t1 20.826
R24355 a_4972_4148.n2 a_4972_4148.n1 20.689
R24356 a_4877_4133.n0 a_4877_4133.t2 362.857
R24357 a_4877_4133.t4 a_4877_4133.t3 337.399
R24358 a_4877_4133.t3 a_4877_4133.t5 298.839
R24359 a_4877_4133.n0 a_4877_4133.t4 280.405
R24360 a_4877_4133.n1 a_4877_4133.t0 200
R24361 a_4877_4133.n1 a_4877_4133.n0 172.311
R24362 a_4877_4133.n2 a_4877_4133.n1 24
R24363 a_4877_4133.n1 a_4877_4133.t1 21.212
R24364 a_6602_n1068.n0 a_6602_n1068.t0 362.857
R24365 a_6602_n1068.t4 a_6602_n1068.t5 337.399
R24366 a_6602_n1068.t5 a_6602_n1068.t3 298.839
R24367 a_6602_n1068.n0 a_6602_n1068.t4 280.405
R24368 a_6602_n1068.n1 a_6602_n1068.t2 200
R24369 a_6602_n1068.n1 a_6602_n1068.n0 172.311
R24370 a_6602_n1068.n2 a_6602_n1068.n1 24
R24371 a_6602_n1068.n1 a_6602_n1068.t1 21.212
R24372 a_6615_n1053.t0 a_6615_n1053.t1 242.857
R24373 a_4890_452.t0 a_4890_452.t1 242.857
R24374 a_8997_4148.n0 a_8997_4148.t1 358.166
R24375 a_8997_4148.t4 a_8997_4148.t5 337.399
R24376 a_8997_4148.t5 a_8997_4148.t3 285.986
R24377 a_8997_4148.n0 a_8997_4148.t4 282.573
R24378 a_8997_4148.n1 a_8997_4148.t2 202.857
R24379 a_8997_4148.n1 a_8997_4148.n0 173.817
R24380 a_8997_4148.n1 a_8997_4148.t0 20.826
R24381 a_8997_4148.n2 a_8997_4148.n1 20.689
R24382 a_9367_4148.t0 a_9367_4148.t1 242.857
R24383 a_7642_693.t0 a_7642_693.t1 242.857
R24384 a_3231_n4116.t0 a_3231_n4116.t1 42.707
R24385 a_3740_1216.t0 a_3740_1216.t1 242.857
R24386 a_8902_4430.n0 a_8902_4430.t0 362.857
R24387 a_8902_4430.t5 a_8902_4430.t4 337.399
R24388 a_8902_4430.t4 a_8902_4430.t3 298.839
R24389 a_8902_4430.n0 a_8902_4430.t5 280.405
R24390 a_8902_4430.n1 a_8902_4430.t2 200
R24391 a_8902_4430.n1 a_8902_4430.n0 172.311
R24392 a_8902_4430.n2 a_8902_4430.n1 24
R24393 a_8902_4430.n1 a_8902_4430.t1 21.212
R24394 a_3617_3907.t0 a_3617_3907.t1 242.857
R24395 a_10327_n7825.t0 a_10327_n7825.t1 42.705
R24396 a_4767_n1053.t0 a_4767_n1053.t1 242.857
R24397 a_7959_n6849.t1 a_7959_n6849.t0 42.707
R24398 a_10327_n6849.t1 a_10327_n6849.t0 42.707
R24399 a_4315_4686.t0 a_4315_4686.t1 242.857
R24400 a_4302_1442.n0 a_4302_1442.t1 362.857
R24401 a_4302_1442.t3 a_4302_1442.t5 337.399
R24402 a_4302_1442.t5 a_4302_1442.t4 298.839
R24403 a_4302_1442.n0 a_4302_1442.t3 280.405
R24404 a_4302_1442.n1 a_4302_1442.t0 200
R24405 a_4302_1442.n1 a_4302_1442.n0 172.311
R24406 a_4302_1442.n2 a_4302_1442.n1 24
R24407 a_4302_1442.n1 a_4302_1442.t2 21.212
R24408 a_8340_1457.t0 a_8340_1457.t1 242.857
R24409 a_1317_693.t0 a_1317_693.t1 242.857
R24410 a_9475_n5338.n0 a_9475_n5338.t0 63.08
R24411 a_9475_n5338.t1 a_9475_n5338.n0 41.303
R24412 a_9475_n5338.n0 a_9475_n5338.t2 2.251
R24413 a_290_3907.t0 a_290_3907.t1 242.857
R24414 a_865_1457.t0 a_865_1457.t1 242.857
R24415 a_3042_211.t0 a_3042_211.t1 242.857
R24416 a_4192_3907.t0 a_4192_3907.t1 242.857
R24417 a_3617_3425.t0 a_3617_3425.t1 242.857
R24418 a_4397_1457.n0 a_4397_1457.t1 358.166
R24419 a_4397_1457.t4 a_4397_1457.t5 337.399
R24420 a_4397_1457.t5 a_4397_1457.t3 285.986
R24421 a_4397_1457.n0 a_4397_1457.t4 282.573
R24422 a_4397_1457.n1 a_4397_1457.t2 202.857
R24423 a_4397_1457.n1 a_4397_1457.n0 173.817
R24424 a_4397_1457.n1 a_4397_1457.t0 20.826
R24425 a_4397_1457.n2 a_4397_1457.n1 20.689
R24426 a_4767_1457.t0 a_4767_1457.t1 242.857
R24427 a_7994_n5293.n0 a_7994_n5293.t0 65.063
R24428 a_7994_n5293.n0 a_7994_n5293.t2 42.011
R24429 a_7994_n5293.t1 a_7994_n5293.n0 2.113
R24430 a_3740_4445.t0 a_3740_4445.t1 242.857
R24431 a_3563_n7203.n0 a_3563_n7203.t0 63.08
R24432 a_3563_n7203.t1 a_3563_n7203.n0 41.306
R24433 a_3563_n7203.n0 a_3563_n7203.t2 2.251
R24434 a_2015_n512.t0 a_2015_n512.t1 242.857
R24435 a_14131_n6847.t1 a_14131_n6847.t0 336.812
R24436 a_13934_n7203.n0 a_13934_n7203.t1 63.08
R24437 a_13934_n7203.t0 a_13934_n7203.n0 41.306
R24438 a_13934_n7203.n0 a_13934_n7203.t2 2.251
R24439 a_7642_3907.t0 a_7642_3907.t1 242.857
R24440 a_7752_3651.n0 a_7752_3651.t0 362.857
R24441 a_7752_3651.t3 a_7752_3651.t4 337.399
R24442 a_7752_3651.t4 a_7752_3651.t5 298.839
R24443 a_7752_3651.n0 a_7752_3651.t3 280.405
R24444 a_7752_3651.n1 a_7752_3651.t2 200
R24445 a_7752_3651.n1 a_7752_3651.n0 172.311
R24446 a_7752_3651.n2 a_7752_3651.n1 24
R24447 a_7752_3651.n1 a_7752_3651.t1 21.212
R24448 a_290_3425.t0 a_290_3425.t1 242.857
R24449 a_1440_3184.t0 a_1440_3184.t1 242.857
R24450 a_5342_975.t0 a_5342_975.t1 242.857
R24451 a_10856_n8026.t1 a_10856_n8026.t0 336.814
R24452 a_10797_n8071.t0 a_10797_n8071.t1 68.74
R24453 a_5465_n271.t0 a_5465_n271.t1 242.857
R24454 a_4192_3425.t0 a_4192_3425.t1 242.857
R24455 a_8997_1698.n0 a_8997_1698.t2 358.166
R24456 a_8997_1698.t4 a_8997_1698.t5 337.399
R24457 a_8997_1698.t5 a_8997_1698.t3 285.986
R24458 a_8997_1698.n0 a_8997_1698.t4 282.573
R24459 a_8997_1698.n1 a_8997_1698.t0 202.857
R24460 a_8997_1698.n1 a_8997_1698.n0 173.817
R24461 a_8997_1698.n1 a_8997_1698.t1 20.826
R24462 a_8997_1698.n2 a_8997_1698.n1 20.689
R24463 a_9367_1698.t0 a_9367_1698.t1 242.857
R24464 a_4302_4671.n0 a_4302_4671.t1 362.857
R24465 a_4302_4671.t3 a_4302_4671.t5 337.399
R24466 a_4302_4671.t5 a_4302_4671.t4 298.839
R24467 a_4302_4671.n0 a_4302_4671.t3 280.405
R24468 a_4302_4671.n1 a_4302_4671.t0 200
R24469 a_4302_4671.n1 a_4302_4671.n0 172.311
R24470 a_4302_4671.n2 a_4302_4671.n1 24
R24471 a_4302_4671.n1 a_4302_4671.t2 21.212
R24472 a_7847_3666.n0 a_7847_3666.t1 358.166
R24473 a_7847_3666.t4 a_7847_3666.t5 337.399
R24474 a_7847_3666.t5 a_7847_3666.t3 285.986
R24475 a_7847_3666.n0 a_7847_3666.t4 282.573
R24476 a_7847_3666.n1 a_7847_3666.t2 202.857
R24477 a_7847_3666.n1 a_7847_3666.n0 173.817
R24478 a_7847_3666.n1 a_7847_3666.t0 20.826
R24479 a_7847_3666.n2 a_7847_3666.n1 20.689
R24480 a_8217_3666.t0 a_8217_3666.t1 242.857
R24481 a_2015_2943.t0 a_2015_2943.t1 242.857
R24482 a_8340_4686.t0 a_8340_4686.t1 242.857
R24483 a_5342_n30.t0 a_5342_n30.t1 242.857
R24484 a_3350_n2132.n0 a_3350_n2132.t2 489.336
R24485 a_3350_n2132.n0 a_3350_n2132.t1 243.258
R24486 a_3350_n2132.t0 a_3350_n2132.n0 214.415
R24487 a_865_4686.t0 a_865_4686.t1 242.857
R24488 Din[3].n0 Din[3].t0 215.292
R24489 Din[3].n0 Din[3].t1 187.376
R24490 Din[3] Din[3].n0 84.903
R24491 a_4397_4686.n0 a_4397_4686.t1 358.166
R24492 a_4397_4686.t4 a_4397_4686.t5 337.399
R24493 a_4397_4686.t5 a_4397_4686.t3 285.986
R24494 a_4397_4686.n0 a_4397_4686.t4 282.573
R24495 a_4397_4686.n1 a_4397_4686.t2 202.857
R24496 a_4397_4686.n1 a_4397_4686.n0 173.817
R24497 a_4397_4686.n1 a_4397_4686.t0 20.826
R24498 a_4397_4686.n2 a_4397_4686.n1 20.689
R24499 a_4767_4686.t0 a_4767_4686.t1 242.857
R24500 a_9613_n5338.t0 a_9613_n5338.t1 68.74
R24501 a_8902_2406.n0 a_8902_2406.t0 362.857
R24502 a_8902_2406.t5 a_8902_2406.t4 337.399
R24503 a_8902_2406.t4 a_8902_2406.t3 298.839
R24504 a_8902_2406.n0 a_8902_2406.t5 280.405
R24505 a_8902_2406.n1 a_8902_2406.t2 200
R24506 a_8902_2406.n1 a_8902_2406.n0 172.311
R24507 a_8902_2406.n2 a_8902_2406.n1 24
R24508 a_8902_2406.n1 a_8902_2406.t1 21.212
R24509 a_8915_n271.t0 a_8915_n271.t1 242.857
R24510 a_8792_1457.t0 a_8792_1457.t1 242.857
R24511 a_7642_3425.t0 a_7642_3425.t1 242.857
R24512 a_3617_n812.t0 a_3617_n812.t1 242.857
R24513 a_13230_n8026.t1 a_13230_n8026.t0 336.814
R24514 a_13171_n8071.t0 a_13171_n8071.t1 68.74
R24515 a_6225_n2132.n0 a_6225_n2132.t2 489.336
R24516 a_6225_n2132.n0 a_6225_n2132.t1 243.258
R24517 a_6225_n2132.t0 a_6225_n2132.n0 214.415
R24518 a_13602_n4116.t0 a_13602_n4116.t1 42.707
R24519 a_8997_1216.n0 a_8997_1216.t2 358.166
R24520 a_8997_1216.t4 a_8997_1216.t5 337.399
R24521 a_8997_1216.t5 a_8997_1216.t3 285.986
R24522 a_8997_1216.n0 a_8997_1216.t4 282.573
R24523 a_8997_1216.n1 a_8997_1216.t0 202.857
R24524 a_8997_1216.n1 a_8997_1216.n0 173.817
R24525 a_8997_1216.n1 a_8997_1216.t1 20.826
R24526 a_8997_1216.n2 a_8997_1216.n1 20.689
R24527 a_9367_1216.t0 a_9367_1216.t1 242.857
R24528 a_865_211.t0 a_865_211.t1 242.857
R24529 a_6040_n512.t0 a_6040_n512.t1 242.857
R24530 a_18_n8071.n0 a_18_n8071.t0 63.08
R24531 a_18_n8071.n0 a_18_n8071.t2 41.307
R24532 a_18_n8071.t1 a_18_n8071.n0 2.251
R24533 a_9367_211.t0 a_9367_211.t1 242.857
R24534 a_4500_n2132.n0 a_4500_n2132.t2 489.336
R24535 a_4500_n2132.n0 a_4500_n2132.t1 243.258
R24536 a_4500_n2132.t0 a_4500_n2132.n0 214.415
R24537 a_4315_2662.t0 a_4315_2662.t1 242.857
R24538 a_2467_n512.t0 a_2467_n512.t1 242.857
R24539 Din[5].n0 Din[5].t0 215.292
R24540 Din[5].n0 Din[5].t1 187.376
R24541 Din[5] Din[5].n0 84.938
R24542 a_2590_4148.t0 a_2590_4148.t1 242.857
R24543 a_290_n812.t0 a_290_n812.t1 242.857
R24544 a_4192_n812.t0 a_4192_n812.t1 242.857
R24545 a_1892_3184.t0 a_1892_3184.t1 242.857
R24546 a_3563_n4470.n0 a_3563_n4470.t0 63.08
R24547 a_3563_n4470.n0 a_3563_n4470.t2 41.305
R24548 a_3563_n4470.t1 a_3563_n4470.n0 2.251
R24549 a_3493_n4483.n0 a_3493_n4483.t3 1464.36
R24550 a_3493_n4483.n0 a_3493_n4483.t4 713.588
R24551 a_3493_n4483.n1 a_3493_n4483.t0 374.998
R24552 a_3493_n4483.n1 a_3493_n4483.t1 273.351
R24553 a_3493_n4483.n2 a_3493_n4483.n0 143.764
R24554 a_3493_n4483.t2 a_3493_n4483.n2 78.209
R24555 a_3493_n4483.n2 a_3493_n4483.n1 4.517
R24556 a_7375_n2132.n0 a_7375_n2132.t2 489.336
R24557 a_7375_n2132.n0 a_7375_n2132.t1 243.258
R24558 a_7375_n2132.t0 a_7375_n2132.n0 214.415
R24559 a_8028_n1770.t0 a_8028_n1770.t1 256.142
R24560 a_3740_2421.t0 a_3740_2421.t1 242.857
R24561 ADC10_OUT[1].n0 ADC10_OUT[1].t4 1355.37
R24562 ADC10_OUT[1].n0 ADC10_OUT[1].t3 820.859
R24563 ADC10_OUT[1].n3 ADC10_OUT[1].t0 330.644
R24564 ADC10_OUT[1].n2 ADC10_OUT[1].t1 266.644
R24565 ADC10_OUT[1].n1 ADC10_OUT[1].n0 149.035
R24566 ADC10_OUT[1].n3 ADC10_OUT[1].n2 53.458
R24567 ADC10_OUT[1] ADC10_OUT[1].n3 46.008
R24568 ADC10_OUT[1].n1 ADC10_OUT[1].t2 45.968
R24569 ADC10_OUT[1].n2 ADC10_OUT[1].n1 17.317
R24570 a_6040_2943.t0 a_6040_2943.t1 242.857
R24571 a_n3298_n6847.t1 a_n3298_n6847.t0 336.812
R24572 a_14131_n4114.t1 a_14131_n4114.t0 336.812
R24573 a_13934_n4470.n0 a_13934_n4470.t0 63.08
R24574 a_13934_n4470.n0 a_13934_n4470.t2 41.305
R24575 a_13934_n4470.t1 a_13934_n4470.n0 2.251
R24576 a_12963_n7216.n0 a_12963_n7216.t4 1464.36
R24577 a_12963_n7216.n0 a_12963_n7216.t3 713.588
R24578 a_12963_n7216.n1 a_12963_n7216.t0 374.998
R24579 a_12963_n7216.n1 a_12963_n7216.t2 273.351
R24580 a_12963_n7216.n2 a_12963_n7216.n0 143.764
R24581 a_12963_n7216.t1 a_12963_n7216.n2 78.209
R24582 a_12963_n7216.n2 a_12963_n7216.n1 4.517
R24583 a_6615_452.t0 a_6615_452.t1 242.857
R24584 a_5917_n512.t0 a_5917_n512.t1 242.857
R24585 a_8792_4686.t0 a_8792_4686.t1 242.857
R24586 a_2097_2943.n0 a_2097_2943.t2 358.166
R24587 a_2097_2943.t4 a_2097_2943.t5 337.399
R24588 a_2097_2943.t5 a_2097_2943.t3 285.986
R24589 a_2097_2943.n0 a_2097_2943.t4 282.573
R24590 a_2097_2943.n1 a_2097_2943.t0 202.857
R24591 a_2097_2943.n1 a_2097_2943.n0 173.817
R24592 a_2097_2943.n1 a_2097_2943.t1 20.826
R24593 a_2097_2943.n2 a_2097_2943.n1 20.689
R24594 a_2467_2943.t0 a_2467_2943.t1 242.857
R24595 a_1317_2180.t0 a_1317_2180.t1 242.857
R24596 a_7642_n812.t0 a_7642_n812.t1 242.857
R24597 a_8997_4445.n0 a_8997_4445.t2 358.166
R24598 a_8997_4445.t4 a_8997_4445.t5 337.399
R24599 a_8997_4445.t5 a_8997_4445.t3 285.986
R24600 a_8997_4445.n0 a_8997_4445.t4 282.573
R24601 a_8997_4445.n1 a_8997_4445.t0 202.857
R24602 a_8997_4445.n1 a_8997_4445.n0 173.817
R24603 a_8997_4445.n1 a_8997_4445.t1 20.826
R24604 a_8997_4445.n2 a_8997_4445.n1 20.689
R24605 a_9367_4445.t0 a_9367_4445.t1 242.857
R24606 a_7765_1939.t0 a_7765_1939.t1 242.857
R24607 a_9178_n1770.n0 a_9178_n1770.t1 160.619
R24608 a_9178_n1770.t0 a_9178_n1770.n0 151.153
R24609 a_5917_2943.t0 a_5917_2943.t1 242.857
R24610 a_4302_2647.n0 a_4302_2647.t1 362.857
R24611 a_4302_2647.t3 a_4302_2647.t5 337.399
R24612 a_4302_2647.t5 a_4302_2647.t4 298.839
R24613 a_4302_2647.n0 a_4302_2647.t3 280.405
R24614 a_4302_2647.n1 a_4302_2647.t0 200
R24615 a_4302_2647.n1 a_4302_2647.n0 172.311
R24616 a_4302_2647.n2 a_4302_2647.n1 24
R24617 a_4302_2647.n1 a_4302_2647.t2 21.212
R24618 a_5768_n2086.t0 a_5768_n2086.t1 34.8
R24619 a_8340_2662.t0 a_8340_2662.t1 242.857
R24620 a_4767_211.t0 a_4767_211.t1 242.857
R24621 a_2519_n4470.t0 a_2519_n4470.t1 68.741
R24622 a_1440_n1053.t0 a_1440_n1053.t1 242.857
R24623 a_6492_n512.t0 a_6492_n512.t1 242.857
R24624 a_865_2662.t0 a_865_2662.t1 242.857
R24625 a_4397_2662.n0 a_4397_2662.t1 358.166
R24626 a_4397_2662.t4 a_4397_2662.t5 337.399
R24627 a_4397_2662.t5 a_4397_2662.t3 285.986
R24628 a_4397_2662.n0 a_4397_2662.t4 282.573
R24629 a_4397_2662.n1 a_4397_2662.t2 202.857
R24630 a_4397_2662.n1 a_4397_2662.n0 173.817
R24631 a_4397_2662.n1 a_4397_2662.t0 20.826
R24632 a_4397_2662.n2 a_4397_2662.n1 20.689
R24633 a_4767_2662.t0 a_4767_2662.t1 242.857
R24634 a_7067_3184.t0 a_7067_3184.t1 242.857
R24635 a_10797_n5338.t0 a_10797_n5338.t1 68.74
R24636 a_742_693.t0 a_742_693.t1 242.857
R24637 a_n2415_n4483.n0 a_n2415_n4483.t3 1464.36
R24638 a_n2415_n4483.n0 a_n2415_n4483.t4 713.588
R24639 a_n2415_n4483.n1 a_n2415_n4483.t0 374.998
R24640 a_n2415_n4483.n1 a_n2415_n4483.t2 273.351
R24641 a_n2415_n4483.n2 a_n2415_n4483.n0 143.764
R24642 a_n2415_n4483.t1 a_n2415_n4483.n2 78.209
R24643 a_n2415_n4483.n2 a_n2415_n4483.n1 4.517
R24644 a_8643_n2086.t0 a_8643_n2086.t1 34.8
R24645 a_6492_452.t0 a_6492_452.t1 242.857
R24646 a_12043_n6847.t1 a_12043_n6847.t0 336.812
R24647 a_6685_n1770.n0 a_6685_n1770.t2 325.682
R24648 a_6685_n1770.t0 a_6685_n1770.n0 322.293
R24649 a_6685_n1770.n0 a_6685_n1770.t1 73.623
R24650 a_2015_3907.t0 a_2015_3907.t1 242.857
R24651 a_6492_2943.t0 a_6492_2943.t1 242.857
R24652 a_6918_n2086.t0 a_6918_n2086.t1 34.8
R24653 a_3165_n1053.t0 a_3165_n1053.t1 242.857
R24654 a_1396_n6847.t1 a_1396_n6847.t0 336.812
R24655 a_1199_n7203.n0 a_1199_n7203.t0 63.08
R24656 a_1199_n7203.n0 a_1199_n7203.t2 41.305
R24657 a_1199_n7203.t1 a_1199_n7203.n0 2.251
R24658 a_5342_2180.t0 a_5342_2180.t1 242.857
R24659 a_2590_1698.t0 a_2590_1698.t1 242.857
R24660 a_n3298_n4114.t1 a_n3298_n4114.t0 336.812
R24661 a_1440_3666.t0 a_1440_3666.t1 242.857
R24662 a_13171_n5338.t0 a_13171_n5338.t1 68.74
R24663 a_3165_1457.t0 a_3165_1457.t1 242.857
R24664 a_2015_3425.t0 a_2015_3425.t1 242.857
R24665 Din[15].n0 Din[15].t0 215.292
R24666 Din[15].n0 Din[15].t1 187.376
R24667 Din[15] Din[15].n0 84.947
R24668 a_8792_2662.t0 a_8792_2662.t1 242.857
R24669 a_5465_975.t0 a_5465_975.t1 242.857
R24670 a_11514_n4116.t0 a_11514_n4116.t1 42.707
R24671 a_2590_1216.t0 a_2590_1216.t1 242.857
R24672 a_8997_2421.n0 a_8997_2421.t2 358.166
R24673 a_8997_2421.t4 a_8997_2421.t5 337.399
R24674 a_8997_2421.t5 a_8997_2421.t3 285.986
R24675 a_8997_2421.n0 a_8997_2421.t4 282.573
R24676 a_8997_2421.n1 a_8997_2421.t0 202.857
R24677 a_8997_2421.n1 a_8997_2421.n0 173.817
R24678 a_8997_2421.n1 a_8997_2421.t1 20.826
R24679 a_8997_2421.n2 a_8997_2421.n1 20.689
R24680 a_9367_2421.t0 a_9367_2421.t1 242.857
R24681 a_1892_452.t0 a_1892_452.t1 242.857
R24682 a_13864_n4483.n0 a_13864_n4483.t3 1464.36
R24683 a_13864_n4483.n0 a_13864_n4483.t4 713.588
R24684 a_13864_n4483.n1 a_13864_n4483.t0 374.998
R24685 a_13864_n4483.n1 a_13864_n4483.t2 273.351
R24686 a_13864_n4483.n2 a_13864_n4483.n0 143.764
R24687 a_13864_n4483.t1 a_13864_n4483.n2 78.209
R24688 a_13864_n4483.n2 a_13864_n4483.n1 4.517
R24689 a_2002_3892.n0 a_2002_3892.t1 362.857
R24690 a_2002_3892.t3 a_2002_3892.t5 337.399
R24691 a_2002_3892.t5 a_2002_3892.t4 298.839
R24692 a_2002_3892.n0 a_2002_3892.t3 280.405
R24693 a_2002_3892.n1 a_2002_3892.t0 200
R24694 a_2002_3892.n1 a_2002_3892.n0 172.311
R24695 a_2002_3892.n2 a_2002_3892.n1 24
R24696 a_2002_3892.n1 a_2002_3892.t2 21.212
R24697 a_6040_3907.t0 a_6040_3907.t1 242.857
R24698 a_4302_2928.n0 a_4302_2928.t1 362.857
R24699 a_4302_2928.t3 a_4302_2928.t5 337.399
R24700 a_4302_2928.t5 a_4302_2928.t4 298.839
R24701 a_4302_2928.n0 a_4302_2928.t3 280.405
R24702 a_4302_2928.n1 a_4302_2928.t0 200
R24703 a_4302_2928.n1 a_4302_2928.n0 172.311
R24704 a_4302_2928.n2 a_4302_2928.n1 24
R24705 a_4302_2928.n1 a_4302_2928.t2 21.212
R24706 a_6615_1457.t0 a_6615_1457.t1 242.857
R24707 a_4883_n4470.t0 a_4883_n4470.t1 68.741
R24708 a_n279_n8026.n0 a_n279_n8026.t0 65.063
R24709 a_n279_n8026.n0 a_n279_n8026.t2 42.011
R24710 a_n279_n8026.t1 a_n279_n8026.n0 2.113
R24711 a_n3495_n5338.n0 a_n3495_n5338.t0 63.08
R24712 a_n3495_n5338.n0 a_n3495_n5338.t2 41.307
R24713 a_n3495_n5338.t1 a_n3495_n5338.n0 2.251
R24714 a_n3357_n5338.t0 a_n3357_n5338.t1 68.74
R24715 a_2097_3907.n0 a_2097_3907.t1 358.166
R24716 a_2097_3907.t4 a_2097_3907.t5 337.399
R24717 a_2097_3907.t5 a_2097_3907.t3 285.986
R24718 a_2097_3907.n0 a_2097_3907.t4 282.573
R24719 a_2097_3907.n1 a_2097_3907.t2 202.857
R24720 a_2097_3907.n1 a_2097_3907.n0 173.817
R24721 a_2097_3907.n1 a_2097_3907.t0 20.826
R24722 a_2097_3907.n2 a_2097_3907.n1 20.689
R24723 a_2467_3907.t0 a_2467_3907.t1 242.857
R24724 a_742_4148.t0 a_742_4148.t1 242.857
R24725 a_9475_n8071.n0 a_9475_n8071.t0 63.08
R24726 a_9475_n8071.t1 a_9475_n8071.n0 41.303
R24727 a_9475_n8071.n0 a_9475_n8071.t2 2.251
R24728 a_7247_n4470.t0 a_7247_n4470.t1 68.741
R24729 a_n314_n7825.t0 a_n314_n7825.t1 42.705
R24730 a_12043_n4114.t1 a_12043_n4114.t0 336.812
R24731 a_3165_4686.t0 a_3165_4686.t1 242.857
R24732 a_1892_3666.t0 a_1892_3666.t1 242.857
R24733 a_2002_3410.n0 a_2002_3410.t1 362.857
R24734 a_2002_3410.t3 a_2002_3410.t5 337.399
R24735 a_2002_3410.t5 a_2002_3410.t4 298.839
R24736 a_2002_3410.n0 a_2002_3410.t3 280.405
R24737 a_2002_3410.n1 a_2002_3410.t0 200
R24738 a_2002_3410.n1 a_2002_3410.n0 172.311
R24739 a_2002_3410.n2 a_2002_3410.n1 24
R24740 a_2002_3410.n1 a_2002_3410.t2 21.212
R24741 a_6040_3425.t0 a_6040_3425.t1 242.857
R24742 a_7190_1457.t0 a_7190_1457.t1 242.857
R24743 a_1396_n4114.t1 a_1396_n4114.t0 336.812
R24744 a_1199_n4470.n0 a_1199_n4470.t0 63.08
R24745 a_1199_n4470.n0 a_1199_n4470.t2 41.305
R24746 a_1199_n4470.t1 a_1199_n4470.n0 2.251
R24747 a_2015_n812.t0 a_2015_n812.t1 242.857
R24748 a_5917_3907.t0 a_5917_3907.t1 242.857
R24749 a_2097_3425.n0 a_2097_3425.t2 358.166
R24750 a_2097_3425.t4 a_2097_3425.t5 337.399
R24751 a_2097_3425.t5 a_2097_3425.t3 285.986
R24752 a_2097_3425.n0 a_2097_3425.t4 282.573
R24753 a_2097_3425.n1 a_2097_3425.t0 202.857
R24754 a_2097_3425.n1 a_2097_3425.n0 173.817
R24755 a_2097_3425.n1 a_2097_3425.t1 20.826
R24756 a_2097_3425.n2 a_2097_3425.n1 20.689
R24757 a_2467_3425.t0 a_2467_3425.t1 242.857
R24758 a_3760_n6847.t1 a_3760_n6847.t0 336.812
R24759 a_2590_4445.t0 a_2590_4445.t1 242.857
R24760 a_6124_n6847.t1 a_6124_n6847.t0 336.812
R24761 a_5927_n7203.n0 a_5927_n7203.t1 63.08
R24762 a_5927_n7203.t0 a_5927_n7203.n0 41.306
R24763 a_5927_n7203.n0 a_5927_n7203.t2 2.251
R24764 a_8902_3169.n0 a_8902_3169.t1 362.857
R24765 a_8902_3169.t5 a_8902_3169.t4 337.399
R24766 a_8902_3169.t4 a_8902_3169.t3 298.839
R24767 a_8902_3169.n0 a_8902_3169.t5 280.405
R24768 a_8902_3169.n1 a_8902_3169.t0 200
R24769 a_8902_3169.n1 a_8902_3169.n0 172.311
R24770 a_8902_3169.n2 a_8902_3169.n1 24
R24771 a_8902_3169.n1 a_8902_3169.t2 21.212
R24772 a_6615_4686.t0 a_6615_4686.t1 242.857
R24773 a_6602_1442.n0 a_6602_1442.t1 362.857
R24774 a_6602_1442.t3 a_6602_1442.t5 337.399
R24775 a_6602_1442.t5 a_6602_1442.t4 298.839
R24776 a_6602_1442.n0 a_6602_1442.t3 280.405
R24777 a_6602_1442.n1 a_6602_1442.t0 200
R24778 a_6602_1442.n1 a_6602_1442.n0 172.311
R24779 a_6602_1442.n2 a_6602_1442.n1 24
R24780 a_6602_1442.n1 a_6602_1442.t2 21.212
R24781 a_9143_n5092.t0 a_9143_n5092.t1 42.705
R24782 a_9178_n5293.n0 a_9178_n5293.t0 65.064
R24783 a_9178_n5293.t1 a_9178_n5293.n0 42.011
R24784 a_9178_n5293.n0 a_9178_n5293.t2 2.113
R24785 a_n279_n5293.n0 a_n279_n5293.t0 65.063
R24786 a_n279_n5293.n0 a_n279_n5293.t2 42.011
R24787 a_n279_n5293.t1 a_n279_n5293.n0 2.113
R24788 a_6492_3907.t0 a_6492_3907.t1 242.857
R24789 a_5917_3425.t0 a_5917_3425.t1 242.857
R24790 a_5465_693.t0 a_5465_693.t1 242.857
R24791 a_3266_n6503.n0 a_3266_n6503.t0 65.064
R24792 a_3266_n6503.n0 a_3266_n6503.t2 42.011
R24793 a_3266_n6503.t1 a_3266_n6503.n0 2.113
R24794 a_7190_211.t0 a_7190_211.t1 242.857
R24795 a_7067_3666.t0 a_7067_3666.t1 242.857
R24796 a_7752_1924.n0 a_7752_1924.t0 362.857
R24797 a_7752_1924.t3 a_7752_1924.t4 337.399
R24798 a_7752_1924.t4 a_7752_1924.t5 298.839
R24799 a_7752_1924.n0 a_7752_1924.t3 280.405
R24800 a_7752_1924.n1 a_7752_1924.t2 200
R24801 a_7752_1924.n1 a_7752_1924.n0 172.311
R24802 a_7752_1924.n2 a_7752_1924.n1 24
R24803 a_7752_1924.n1 a_7752_1924.t1 21.212
R24804 a_n1460_n8026.n0 a_n1460_n8026.t0 65.063
R24805 a_n1460_n8026.n0 a_n1460_n8026.t2 42.011
R24806 a_n1460_n8026.t1 a_n1460_n8026.n0 2.113
R24807 a_4315_n512.t0 a_4315_n512.t1 242.857
R24808 a_7190_4686.t0 a_7190_4686.t1 242.857
R24809 a_1128_n1770.t0 a_1128_n1770.t1 256.142
R24810 Din[0].n0 Din[0].t0 215.292
R24811 Din[0].n0 Din[0].t1 187.376
R24812 Din[0] Din[0].n0 85.063
R24813 a_6040_n812.t0 a_6040_n812.t1 242.857
R24814 a_6697_n1053.n0 a_6697_n1053.t1 358.166
R24815 a_6697_n1053.t3 a_6697_n1053.t4 337.399
R24816 a_6697_n1053.t4 a_6697_n1053.t5 285.986
R24817 a_6697_n1053.n0 a_6697_n1053.t3 282.573
R24818 a_6697_n1053.n1 a_6697_n1053.t2 202.857
R24819 a_6697_n1053.n1 a_6697_n1053.n0 173.817
R24820 a_6697_n1053.n1 a_6697_n1053.t0 20.826
R24821 a_6697_n1053.n2 a_6697_n1053.n1 20.689
R24822 a_3740_3184.t0 a_3740_3184.t1 242.857
R24823 a_7765_n271.t0 a_7765_n271.t1 242.857
R24824 a_5595_n4116.t0 a_5595_n4116.t1 42.707
R24825 a_1892_n30.t0 a_1892_n30.t1 242.857
R24826 a_6492_3425.t0 a_6492_3425.t1 242.857
R24827 a_2467_n812.t0 a_2467_n812.t1 242.857
R24828 a_8217_452.t0 a_8217_452.t1 242.857
R24829 ADC4_OUT[2].n0 ADC4_OUT[2].t4 1354.27
R24830 ADC4_OUT[2].n0 ADC4_OUT[2].t3 821.954
R24831 ADC4_OUT[2].n3 ADC4_OUT[2].t0 347.891
R24832 ADC4_OUT[2].n2 ADC4_OUT[2].t2 266.575
R24833 ADC4_OUT[2].n1 ADC4_OUT[2].n0 149.035
R24834 ADC4_OUT[2].n1 ADC4_OUT[2].t1 46.723
R24835 ADC4_OUT[2] ADC4_OUT[2].n3 37.824
R24836 ADC4_OUT[2].n3 ADC4_OUT[2].n2 36.141
R24837 ADC4_OUT[2].n2 ADC4_OUT[2].n1 17.317
R24838 a_4003_n1770.t0 a_4003_n1770.t1 256.142
R24839 a_6602_4671.n0 a_6602_4671.t1 362.857
R24840 a_6602_4671.t3 a_6602_4671.t5 337.399
R24841 a_6602_4671.t5 a_6602_4671.t4 298.839
R24842 a_6602_4671.n0 a_6602_4671.t3 280.405
R24843 a_6602_4671.n1 a_6602_4671.t0 200
R24844 a_6602_4671.n1 a_6602_4671.n0 172.311
R24845 a_6602_4671.n2 a_6602_4671.n1 24
R24846 a_6602_4671.n1 a_6602_4671.t2 21.212
R24847 a_4315_2943.t0 a_4315_2943.t1 242.857
R24848 a_10659_n8071.n0 a_10659_n8071.t0 63.08
R24849 a_10659_n8071.n0 a_10659_n8071.t2 41.307
R24850 a_10659_n8071.t1 a_10659_n8071.n0 2.251
R24851 a_742_1698.t0 a_742_1698.t1 242.857
R24852 a_5628_n2086.t0 a_5628_n2086.t1 34.8
R24853 a_3165_2662.t0 a_3165_2662.t1 242.857
R24854 a_6697_1457.n0 a_6697_1457.t1 358.166
R24855 a_6697_1457.t3 a_6697_1457.t4 337.399
R24856 a_6697_1457.t4 a_6697_1457.t5 285.986
R24857 a_6697_1457.n0 a_6697_1457.t3 282.573
R24858 a_6697_1457.n1 a_6697_1457.t2 202.857
R24859 a_6697_1457.n1 a_6697_1457.n0 173.817
R24860 a_6697_1457.n1 a_6697_1457.t0 20.826
R24861 a_6697_1457.n2 a_6697_1457.n1 20.689
R24862 a_n966_n5293.t1 a_n966_n5293.t0 336.814
R24863 a_2278_n1770.n0 a_2278_n1770.t1 160.619
R24864 a_2278_n1770.t0 a_2278_n1770.n0 151.153
R24865 a_3760_n4114.t1 a_3760_n4114.t0 336.812
R24866 a_5917_n812.t0 a_5917_n812.t1 242.857
R24867 a_6124_n4114.t1 a_6124_n4114.t0 336.812
R24868 a_5927_n4470.n0 a_5927_n4470.t0 63.08
R24869 a_5927_n4470.n0 a_5927_n4470.t2 41.305
R24870 a_5927_n4470.t1 a_5927_n4470.n0 2.251
R24871 a_2590_211.t0 a_2590_211.t1 242.857
R24872 a_8503_n2086.t0 a_8503_n2086.t1 34.8
R24873 a_2590_2421.t0 a_2590_2421.t1 242.857
R24874 a_8340_n512.t0 a_8340_n512.t1 242.857
R24875 a_742_1216.t0 a_742_1216.t1 242.857
R24876 a_865_n512.t0 a_865_n512.t1 242.857
R24877 a_6615_2662.t0 a_6615_2662.t1 242.857
R24878 a_4767_n512.t0 a_4767_n512.t1 242.857
R24879 a_12701_n7825.t0 a_12701_n7825.t1 42.705
R24880 a_4890_4148.t0 a_4890_4148.t1 242.857
R24881 a_6492_n812.t0 a_6492_n812.t1 242.857
R24882 a_8915_975.t0 a_8915_975.t1 242.857
R24883 a_865_n30.t0 a_865_n30.t1 242.857
R24884 a_12701_n6849.t0 a_12701_n6849.t1 42.707
R24885 a_3617_452.t0 a_3617_452.t1 242.857
R24886 a_8340_2943.t0 a_8340_2943.t1 242.857
R24887 a_6697_4686.n0 a_6697_4686.t1 358.166
R24888 a_6697_4686.t3 a_6697_4686.t4 337.399
R24889 a_6697_4686.t4 a_6697_4686.t5 285.986
R24890 a_6697_4686.n0 a_6697_4686.t3 282.573
R24891 a_6697_4686.n1 a_6697_4686.t2 202.857
R24892 a_6697_4686.n1 a_6697_4686.n0 173.817
R24893 a_6697_4686.n1 a_6697_4686.t0 20.826
R24894 a_6697_4686.n2 a_6697_4686.n1 20.689
R24895 a_865_2943.t0 a_865_2943.t1 242.857
R24896 a_977_n1770.t0 a_977_n1770.n0 182.779
R24897 a_977_n1770.n0 a_977_n1770.t1 111.474
R24898 a_4397_2943.n0 a_4397_2943.t2 358.166
R24899 a_4397_2943.t4 a_4397_2943.t5 337.399
R24900 a_4397_2943.t5 a_4397_2943.t3 285.986
R24901 a_4397_2943.n0 a_4397_2943.t4 282.573
R24902 a_4397_2943.n1 a_4397_2943.t0 202.857
R24903 a_4397_2943.n1 a_4397_2943.n0 173.817
R24904 a_4397_2943.n1 a_4397_2943.t1 20.826
R24905 a_4397_2943.n2 a_4397_2943.n1 20.689
R24906 a_4767_2943.t0 a_4767_2943.t1 242.857
R24907 a_7190_2662.t0 a_7190_2662.t1 242.857
R24908 a_2893_n2086.t0 a_2893_n2086.t1 34.8
R24909 a_3617_2180.t0 a_3617_2180.t1 242.857
R24910 a_4890_n30.t0 a_4890_n30.t1 242.857
R24911 a_7959_n4116.t0 a_7959_n4116.t1 42.707
R24912 a_10327_n4116.t0 a_10327_n4116.t1 42.707
R24913 a_742_4445.t0 a_742_4445.t1 242.857
R24914 a_7847_1939.n0 a_7847_1939.t1 358.166
R24915 a_7847_1939.t4 a_7847_1939.t5 337.399
R24916 a_7847_1939.t5 a_7847_1939.t3 285.986
R24917 a_7847_1939.n0 a_7847_1939.t4 282.573
R24918 a_7847_1939.n1 a_7847_1939.t2 202.857
R24919 a_7847_1939.n1 a_7847_1939.n0 173.817
R24920 a_7847_1939.n1 a_7847_1939.t0 20.826
R24921 a_7847_1939.n2 a_7847_1939.n1 20.689
R24922 a_8902_3651.n0 a_8902_3651.t0 362.857
R24923 a_8902_3651.t5 a_8902_3651.t4 337.399
R24924 a_8902_3651.t4 a_8902_3651.t3 298.839
R24925 a_8902_3651.n0 a_8902_3651.t5 280.405
R24926 a_8902_3651.n1 a_8902_3651.t2 200
R24927 a_8902_3651.n1 a_8902_3651.n0 172.311
R24928 a_8902_3651.n2 a_8902_3651.n1 24
R24929 a_8902_3651.n1 a_8902_3651.t1 21.212
R24930 a_8792_n512.t0 a_8792_n512.t1 242.857
R24931 a_290_2180.t0 a_290_2180.t1 242.857
R24932 a_8792_975.t0 a_8792_975.t1 242.857
R24933 a_3042_4148.t0 a_3042_4148.t1 242.857
R24934 a_8997_3184.n0 a_8997_3184.t2 358.166
R24935 a_8997_3184.t4 a_8997_3184.t5 337.399
R24936 a_8997_3184.t5 a_8997_3184.t3 285.986
R24937 a_8997_3184.n0 a_8997_3184.t4 282.573
R24938 a_8997_3184.n1 a_8997_3184.t0 202.857
R24939 a_8997_3184.n1 a_8997_3184.n0 173.817
R24940 a_8997_3184.n1 a_8997_3184.t1 20.826
R24941 a_8997_3184.n2 a_8997_3184.n1 20.689
R24942 a_9367_3184.t0 a_9367_3184.t1 242.857
R24943 a_4192_2180.t0 a_4192_2180.t1 242.857
R24944 a_4315_3907.t0 a_4315_3907.t1 242.857
R24945 a_8792_2943.t0 a_8792_2943.t1 242.857
R24946 a_2015_975.t0 a_2015_975.t1 242.857
R24947 a_7642_2180.t0 a_7642_2180.t1 242.857
R24948 a_n2148_n8026.t1 a_n2148_n8026.t0 336.814
R24949 a_8915_693.t0 a_8915_693.t1 242.857
R24950 ADC0_OUT[1].n0 ADC0_OUT[1].t4 1355.37
R24951 ADC0_OUT[1].n0 ADC0_OUT[1].t3 820.859
R24952 ADC0_OUT[1].n3 ADC0_OUT[1].t0 350.973
R24953 ADC0_OUT[1].n2 ADC0_OUT[1].t2 266.644
R24954 ADC0_OUT[1].n1 ADC0_OUT[1].n0 149.035
R24955 ADC0_OUT[1].n1 ADC0_OUT[1].t1 45.968
R24956 ADC0_OUT[1] ADC0_OUT[1].n3 45.82
R24957 ADC0_OUT[1].n3 ADC0_OUT[1].n2 33.129
R24958 ADC0_OUT[1].n2 ADC0_OUT[1].n1 17.317
R24959 a_3740_3666.t0 a_3740_3666.t1 242.857
R24960 a_4890_1698.t0 a_4890_1698.t1 242.857
R24961 a_n1495_n7825.t0 a_n1495_n7825.t1 42.705
R24962 a_8217_1939.t0 a_8217_1939.t1 242.857
R24963 a_215_n6847.t1 a_215_n6847.t0 336.812
R24964 a_2467_975.t0 a_2467_975.t1 242.857
R24965 a_4315_3425.t0 a_4315_3425.t1 242.857
R24966 a_5465_1457.t0 a_5465_1457.t1 242.857
R24967 a_4675_n5850.n0 a_4675_n5850.t4 1465.51
R24968 a_4675_n5850.n0 a_4675_n5850.t3 712.44
R24969 a_4675_n5850.n1 a_4675_n5850.t0 375.067
R24970 a_4675_n5850.n1 a_4675_n5850.t1 272.668
R24971 a_4675_n5850.n2 a_4675_n5850.n0 143.764
R24972 a_4675_n5850.t2 a_4675_n5850.n2 78.193
R24973 a_4675_n5850.n2 a_4675_n5850.n1 4.517
R24974 a_n1025_n7203.t0 a_n1025_n7203.t1 68.741
R24975 a_4890_1216.t0 a_4890_1216.t1 242.857
R24976 a_8340_3907.t0 a_8340_3907.t1 242.857
R24977 a_742_2421.t0 a_742_2421.t1 242.857
R24978 a_8915_1457.t0 a_8915_1457.t1 242.857
R24979 a_7067_693.t0 a_7067_693.t1 242.857
R24980 a_290_211.t0 a_290_211.t1 242.857
R24981 a_865_3907.t0 a_865_3907.t1 242.857
R24982 a_4767_3907.t0 a_4767_3907.t1 242.857
R24983 a_8792_693.t0 a_8792_693.t1 242.857
R24984 a_4315_211.t0 a_4315_211.t1 242.857
R24985 a_14131_n5293.t1 a_14131_n5293.t0 336.814
R24986 a_n314_n5092.t0 a_n314_n5092.t1 42.705
R24987 a_3042_1698.t0 a_3042_1698.t1 242.857
R24988 a_7190_n30.t0 a_7190_n30.t1 242.857
R24989 a_5465_4686.t0 a_5465_4686.t1 242.857
R24990 a_8340_3425.t0 a_8340_3425.t1 242.857
R24991 a_6040_452.t0 a_6040_452.t1 242.857
R24992 a_4315_n812.t0 a_4315_n812.t1 242.857
R24993 a_865_3425.t0 a_865_3425.t1 242.857
R24994 a_5917_975.t0 a_5917_975.t1 242.857
R24995 a_4767_3425.t0 a_4767_3425.t1 242.857
R24996 a_4890_4445.t0 a_4890_4445.t1 242.857
R24997 a_475_n2132.n0 a_475_n2132.t2 489.336
R24998 a_475_n2132.n0 a_475_n2132.t1 243.258
R24999 a_475_n2132.t0 a_475_n2132.n0 214.415
R25000 a_215_n4114.t1 a_215_n4114.t0 336.812
R25001 a_8915_4686.t0 a_8915_4686.t1 242.857
R25002 a_3042_1216.t0 a_3042_1216.t1 242.857
R25003 a_3165_n512.t0 a_3165_n512.t1 242.857
R25004 a_2467_693.t0 a_2467_693.t1 242.857
R25005 a_1603_n2086.t0 a_1603_n2086.t1 34.8
R25006 a_8792_3907.t0 a_8792_3907.t1 242.857
R25007 a_4192_211.t0 a_4192_211.t1 242.857
R25008 a_2590_3184.t0 a_2590_3184.t1 242.857
R25009 a_8997_3666.n0 a_8997_3666.t1 358.166
R25010 a_8997_3666.t4 a_8997_3666.t5 337.399
R25011 a_8997_3666.t5 a_8997_3666.t3 285.986
R25012 a_8997_3666.n0 a_8997_3666.t4 282.573
R25013 a_8997_3666.n1 a_8997_3666.t2 202.857
R25014 a_8997_3666.n1 a_8997_3666.n0 173.817
R25015 a_8997_3666.n1 a_8997_3666.t0 20.826
R25016 a_8997_3666.n2 a_8997_3666.n1 20.689
R25017 a_9367_3666.t0 a_9367_3666.t1 242.857
R25018 a_3165_2943.t0 a_3165_2943.t1 242.857
R25019 a_6615_n512.t0 a_6615_n512.t1 242.857
R25020 a_n3298_n5293.t1 a_n3298_n5293.t0 336.814
R25021 a_6615_2943.t0 a_6615_2943.t1 242.857
R25022 a_1440_1939.t0 a_1440_1939.t1 242.857
R25023 a_9672_n6847.t1 a_9672_n6847.t0 336.812
R25024 a_9475_n7203.n0 a_9475_n7203.t1 63.08
R25025 a_9475_n7203.t0 a_9475_n7203.n0 41.306
R25026 a_9475_n7203.n0 a_9475_n7203.t2 2.251
R25027 a_7190_2943.t0 a_7190_2943.t1 242.857
R25028 a_12043_n5293.t1 a_12043_n5293.t0 336.814
R25029 a_11984_n5338.t0 a_11984_n5338.t1 68.74
R25030 a_1396_n5293.t1 a_1396_n5293.t0 336.814
R25031 a_14072_n7203.t0 a_14072_n7203.t1 68.741
R25032 a_1892_1939.t0 a_1892_1939.t1 242.857
R25033 a_7959_n7825.t0 a_7959_n7825.t1 42.705
R25034 a_10856_n6847.t1 a_10856_n6847.t0 336.812
R25035 a_7067_1939.t0 a_7067_1939.t1 242.857
R25036 a_8488_n8026.t1 a_8488_n8026.t0 336.814
R25037 a_8429_n8071.t0 a_8429_n8071.t1 68.74
R25038 a_13230_n6847.t1 a_13230_n6847.t0 336.812
R25039 a_3760_n5293.t1 a_3760_n5293.t0 336.814
R25040 a_6124_n5293.t1 a_6124_n5293.t0 336.814
R25041 a_6777_n5092.t0 a_6777_n5092.t1 42.705
R25042 a_8340_975.t0 a_8340_975.t1 242.857
R25043 a_12701_n4116.t0 a_12701_n4116.t1 42.707
R25044 a_1337_n7203.t0 a_1337_n7203.t1 68.741
R25045 a_3617_n30.t0 a_3617_n30.t1 242.857
R25046 a_4478_n2086.t0 a_4478_n2086.t1 34.8
R25047 a_9367_n30.t0 a_9367_n30.t1 242.857
R25048 a_3701_n7203.t0 a_3701_n7203.t1 68.741
R25049 a_2084_n5293.n0 a_2084_n5293.t0 65.063
R25050 a_2084_n5293.n0 a_2084_n5293.t2 42.011
R25051 a_2084_n5293.t1 a_2084_n5293.n0 2.113
R25052 a_n1025_n4470.t0 a_n1025_n4470.t1 68.741
R25053 a_6065_n7203.t0 a_6065_n7203.t1 68.741
R25054 a_2702_n1770.t0 a_2702_n1770.t1 213.924
R25055 a_1440_n30.t0 a_1440_n30.t1 242.857
R25056 a_3852_n1770.t0 a_3852_n1770.t1 213.924
R25057 a_215_n5293.t1 a_215_n5293.t0 336.814
R25058 a_3165_975.t0 a_3165_975.t1 242.857
R25059 a_14072_n4470.t0 a_14072_n4470.t1 68.741
R25060 a_4448_n5293.n0 a_4448_n5293.t0 65.063
R25061 a_4448_n5293.n0 a_4448_n5293.t2 42.011
R25062 a_4448_n5293.t1 a_4448_n5293.n0 2.113
R25063 ADC5_OUT[1].n0 ADC5_OUT[1].t4 1355.37
R25064 ADC5_OUT[1].n0 ADC5_OUT[1].t3 820.859
R25065 ADC5_OUT[1].n3 ADC5_OUT[1].t0 331.396
R25066 ADC5_OUT[1].n2 ADC5_OUT[1].t1 266.644
R25067 ADC5_OUT[1].n1 ADC5_OUT[1].n0 149.035
R25068 ADC5_OUT[1].n3 ADC5_OUT[1].n2 52.705
R25069 ADC5_OUT[1].n1 ADC5_OUT[1].t2 45.968
R25070 ADC5_OUT[1] ADC5_OUT[1].n3 45.848
R25071 ADC5_OUT[1].n2 ADC5_OUT[1].n1 17.317
R25072 a_8291_n8071.n0 a_8291_n8071.t0 63.08
R25073 a_8291_n8071.t1 a_8291_n8071.n0 41.303
R25074 a_8291_n8071.n0 a_8291_n8071.t2 2.251
R25075 a_156_n7203.t0 a_156_n7203.t1 68.741
R25076 a_9672_n5293.t1 a_9672_n5293.t0 336.814
R25077 a_1337_n4470.t0 a_1337_n4470.t1 68.741
R25078 a_7493_n2086.t0 a_7493_n2086.t1 34.8
R25079 a_10856_n5293.t1 a_10856_n5293.t0 336.814
R25080 a_3701_n4470.t0 a_3701_n4470.t1 68.741
R25081 a_6065_n4470.t0 a_6065_n4470.t1 68.741
R25082 a_13230_n5293.t1 a_13230_n5293.t0 336.814
R25083 a_9613_n7203.t0 a_9613_n7203.t1 68.741
R25084 a_156_n4470.t0 a_156_n4470.t1 68.741
R25085 a_6878_n1770.t0 a_6878_n1770.t1 256.142
C0 a_5632_n6430# Iref0 0.00fF
C1 a_5743_n6391# ADC13_OUT[0] 0.02fF
C2 PRE_CLSA ADC9_OUT[3] 0.10fF
C3 ADC3_OUT[1] ADC3_OUT[2] 3.78fF
C4 a_5632_n6430# VDD 0.98fF
C5 VCLP ADC9_OUT[2] 0.02fF
C6 ADC7_OUT[1] Iref1 0.01fF
C7 ADC9_OUT[0] Iref2 0.01fF
C8 SAEN ADC8_OUT[2] 0.01fF
C9 ADC4_OUT[0] ADC4_OUT[3] 0.03fF
C10 WWL[8] RWLB[9] 0.01fF
C11 RWLB[8] WWL[9] 0.02fF
C12 RWLB[7] WWL[10] 0.01fF
C13 RWL[7] RWL[10] 0.00fF
C14 RWL[8] RWL[9] 0.09fF
C15 VDD SA_OUT[6] 1.34fF
C16 WWL[7] RWLB[10] 0.00fF
C17 VDD ADC7_OUT[2] 1.53fF
C18 a_5632_n6430# ADC10_OUT[1] 0.01fF
C19 a_5743_n6391# Iref1 0.00fF
C20 SAEN ADC13_OUT[3] 0.02fF
C21 ADC8_OUT[1] ADC9_OUT[2] 0.01fF
C22 ADC9_OUT[0] ADC10_OUT[3] 0.00fF
C23 RWL[9] WWL[12] 0.00fF
C24 RWL[10] WWL[11] 0.01fF
C25 RWLB[9] RWLB[11] 0.02fF
C26 WWL[9] RWL[12] 0.01fF
C27 WWL[10] RWL[11] 0.02fF
C28 VDD Din[0] 0.24fF
C29 m1_2243_5034# VDD 0.06fF
C30 ADC13_OUT[0] ADC14_OUT[0] 0.01fF
C31 ADC11_OUT[0] VCLP 0.87fF
C32 a_5743_n6391# ADC10_OUT[2] 0.92fF
C33 ADC0_OUT[2] Iref3 0.01fF
C34 WWL[12] WWL[13] 0.10fF
C35 RWL[12] RWLB[12] 0.08fF
C36 VDD Din[11] 0.26fF
C37 RWL[1] Din[1] 0.01fF
C38 WWLD[0] Din[9] 0.00fF
C39 WWL[1] Din[2] 0.00fF
C40 WWLD[2] Din[7] 0.00fF
C41 WWLD[3] Din[6] 0.00fF
C42 WWLD[1] Din[8] 0.00fF
C43 PRE_SRAM Din[10] 0.01fF
C44 WWL[0] Din[5] 0.00fF
C45 WWL[11] WWL[14] 0.01fF
C46 RWLB[1] Din[0] 0.00fF
C47 RWL[0] Din[4] 0.00fF
C48 RWLB[11] RWL[13] 0.01fF
C49 RWLB[0] Din[3] 0.01fF
C50 RWL[11] RWLB[13] 0.01fF
C51 VCLP ADC14_OUT[1] 0.95fF
C52 ADC15_OUT[0] ADC15_OUT[1] 5.50fF
C53 PRE_CLSA ADC14_OUT[2] 0.09fF
C54 ADC14_OUT[0] Iref1 0.02fF
C55 ADC3_OUT[0] Iref0 0.03fF
C56 ADC5_OUT[0] VCLP 0.89fF
C57 ADC1_OUT[0] ADC1_OUT[1] 5.50fF
C58 PRE_CLSA ADC3_OUT[1] 0.10fF
C59 ADC4_OUT[0] SAEN 0.07fF
C60 WWL[5] Din[1] 0.00fF
C61 RWLB[1] Din[11] 0.01fF
C62 RWLB[4] Din[2] 0.01fF
C63 RWLB[2] Din[8] 0.01fF
C64 VDD ADC3_OUT[0] 2.27fF
C65 WWL[13] RWLB[15] 0.01fF
C66 RWL[2] Din[9] 0.00fF
C67 RWLB[0] Din[14] 0.01fF
C68 RWLB[3] Din[5] 0.01fF
C69 WWL[1] Din[13] 0.00fF
C70 RWL[1] Din[12] 0.00fF
C71 RWL[3] Din[6] 0.00fF
C72 RWL[4] Din[3] 0.01fF
C73 RWL[0] Din[15] 0.00fF
C74 RWL[13] RWL[15] 0.02fF
C75 RWL[5] Din[0] 0.00fF
C76 WWL[2] Din[10] 0.00fF
C77 WWL[14] RWLB[14] 21.69fF
C78 WWL[4] Din[4] 0.00fF
C79 RWLB[13] WWL[15] 0.02fF
C80 WWL[3] Din[7] 0.00fF
C81 ADC12_OUT[0] ADC12_OUT[2] 0.03fF
C82 ADC6_OUT[0] ADC7_OUT[1] 0.00fF
C83 RWLB[15] WWLD[6] 0.00fF
C84 RWL[4] Din[14] 0.00fF
C85 RWLB[5] Din[10] 0.01fF
C86 RWL[5] Din[11] 0.00fF
C87 RWLB[4] Din[13] 0.01fF
C88 WWL[8] Din[3] 0.00fF
C89 WWLD[4] WWLD[5] 0.86fF
C90 WWL[5] Din[12] 0.00fF
C91 RWL[7] Din[5] 0.00fF
C92 RWLB[7] Din[4] 0.01fF
C93 RWL[8] Din[2] 0.00fF
C94 WWL[6] Din[9] 0.00fF
C95 WWL[7] Din[6] 0.00fF
C96 RWL[6] Din[8] 0.00fF
C97 ADC13_OUT[1] ADC14_OUT[2] 0.01fF
C98 RWLB[6] Din[7] 0.01fF
C99 WWL[4] Din[15] 0.00fF
C100 WWL[9] Din[0] 0.00fF
C101 ADC11_OUT[1] Iref2 0.01fF
C102 RWLB[8] Din[1] 0.01fF
C103 VDD ADC11_OUT[3] 1.58fF
C104 m1_1095_5034# PRE_SRAM 0.14fF
C105 RWL[11] Din[4] 0.00fF
C106 RWL[10] Din[7] 0.00fF
C107 RWLB[8] Din[12] 0.01fF
C108 RWLB[10] Din[6] 0.01fF
C109 WWL[11] Din[5] 0.00fF
C110 WWL[9] Din[11] 0.00fF
C111 RWLB[11] Din[3] 0.01fF
C112 RWLB[12] Din[0] 0.00fF
C113 RWLB[7] Din[15] 0.01fF
C114 RWL[12] Din[1] 0.01fF
C115 SA_OUT[0] SA_OUT[2] 0.00fF
C116 ADC10_OUT[1] ADC11_OUT[3] 0.00fF
C117 WWLD[6] SA_OUT[5] 0.03fF
C118 PRE_VLSA SA_OUT[3] 0.17fF
C119 RWL[8] Din[13] 0.00fF
C120 ADC10_OUT[2] ADC11_OUT[2] 0.01fF
C121 WWL[8] Din[14] 0.00fF
C122 RWL[9] Din[10] 0.00fF
C123 RWLB[9] Din[9] 0.01fF
C124 WWLD[5] SA_OUT[6] 0.00fF
C125 WWL[12] Din[2] 0.00fF
C126 WWLD[7] SA_OUT[4] 0.05fF
C127 WWL[10] Din[8] 0.00fF
C128 ADC5_OUT[1] Iref2 0.01fF
C129 ADC7_OUT[0] Iref3 0.01fF
C130 SAEN ADC6_OUT[3] 0.02fF
C131 VCLP ADC7_OUT[3] 1.02fF
C132 ADC2_OUT[1] ADC2_OUT[3] 0.01fF
C133 SAEN ADC12_OUT[1] 0.03fF
C134 VDD ADC5_OUT[3] 1.58fF
C135 a_5632_n6430# ADC8_OUT[2] 0.03fF
C136 WWLD[4] Din[1] 0.00fF
C137 SA_OUT[1] SA_OUT[12] 0.00fF
C138 PRE_VLSA SA_OUT[14] 0.13fF
C139 WWL[15] Din[4] 0.00fF
C140 RWL[14] Din[6] 0.00fF
C141 RWL[15] Din[3] 0.00fF
C142 SA_OUT[0] SA_OUT[13] 0.00fF
C143 RWL[13] Din[9] 0.00fF
C144 SA_OUT[2] SA_OUT[11] 0.01fF
C145 SA_OUT[6] SA_OUT[7] 5.61fF
C146 SA_OUT[5] SA_OUT[8] 0.01fF
C147 RWLB[14] Din[5] 0.01fF
C148 WWL[14] Din[7] 0.00fF
C149 SA_OUT[4] SA_OUT[9] 0.01fF
C150 RWL[12] Din[12] 0.00fF
C151 WWL[13] Din[10] 0.00fF
C152 RWLB[12] Din[11] 0.01fF
C153 RWLB[11] Din[14] 0.01fF
C154 WWLD[5] Din[0] 0.00fF
C155 WWLD[7] SA_OUT[15] 0.02fF
C156 SA_OUT[3] SA_OUT[10] 0.01fF
C157 WWL[12] Din[13] 0.00fF
C158 RWL[11] Din[15] 0.00fF
C159 RWLB[13] Din[8] 0.01fF
C160 RWLB[15] Din[2] 0.01fF
C161 ADC7_OUT[2] ADC8_OUT[2] 0.01fF
C162 ADC7_OUT[1] ADC8_OUT[3] 0.00fF
C163 RWLB[15] Din[13] 0.01fF
C164 SA_OUT[11] SA_OUT[13] 0.01fF
C165 SA_OUT[2] Din[5] 0.01fF
C166 WWLD[5] Din[11] 0.00fF
C167 SA_OUT[3] Din[4] 0.01fF
C168 WWLD[7] Din[9] 0.00fF
C169 WWLD[4] Din[12] 0.00fF
C170 SA_OUT[10] SA_OUT[14] 0.02fF
C171 SA_OUT[0] Din[7] 0.02fF
C172 SA_OUT[9] SA_OUT[15] 0.02fF
C173 WWLD[6] Din[10] 0.00fF
C174 RWL[15] Din[14] 0.00fF
C175 PRE_VLSA Din[8] 0.02fF
C176 SA_OUT[8] WE 0.02fF
C177 SA_OUT[1] Din[6] 0.01fF
C178 WWL[15] Din[15] 0.00fF
C179 SA_OUT[2] PRE_A 0.00fF
C180 SA_OUT[1] EN 0.00fF
C181 SA_OUT[8] Din[10] 0.01fF
C182 SA_OUT[5] Din[13] 0.01fF
C183 Din[0] Din[1] 0.02fF
C184 SA_OUT[7] Din[11] 0.01fF
C185 ADC9_OUT[3] Iref3 0.01fF
C186 WE Din[2] 0.01fF
C187 SA_OUT[6] Din[12] 0.01fF
C188 SA_OUT[9] Din[9] 0.00fF
C189 SA_OUT[4] Din[14] 0.01fF
C190 SA_OUT[3] Din[15] 0.01fF
C191 SAEN ADC0_OUT[1] 0.04fF
C192 ADC0_OUT[0] ADC0_OUT[2] 0.03fF
C193 VCLP ADC1_OUT[1] 0.92fF
C194 PRE_CLSA ADC1_OUT[2] 0.09fF
C195 ADC1_OUT[0] Iref1 0.02fF
C196 VDD Iref0 0.45fF
C197 SA_OUT[14] Din[15] 0.02fF
C198 SA_OUT[12] EN 0.01fF
C199 WE Din[13] 0.01fF
C200 SA_OUT[13] PRE_A 0.01fF
C201 ADC5_OUT[0] ADC6_OUT[2] 0.00fF
C202 Iref0 ADC10_OUT[1] 0.00fF
C203 ADC4_OUT[1] ADC5_OUT[1] 0.01fF
C204 m1_6843_5034# m1_7418_5034# 0.00fF
C205 VDD ADC10_OUT[1] 1.57fF
C206 Din[7] PRE_A 0.00fF
C207 Din[11] Din[12] 0.02fF
C208 Din[6] EN 0.00fF
C209 WWLD[1] RWLB[0] 0.00fF
C210 WWLD[3] WWL[0] 0.10fF
C211 VDD RWLB[1] 2.06fF
C212 WWLD[2] RWL[0] 0.01fF
C213 ADC15_OUT[2] ADC15_OUT[3] 1.31fF
C214 Iref2 ADC14_OUT[3] 0.00fF
C215 ADC14_OUT[2] Iref3 0.01fF
C216 ADC3_OUT[2] Iref2 0.02fF
C217 ADC3_OUT[1] Iref3 0.01fF
C218 ADC1_OUT[2] ADC1_OUT[3] 1.31fF
C219 RWL[0] WWL[3] 0.00fF
C220 RWL[1] WWL[2] 0.01fF
C221 PRE_A PRE_CLSA 0.14fF
C222 WWL[1] RWL[2] 0.02fF
C223 VDD RWL[5] 2.83fF
C224 WWL[0] RWL[3] 0.01fF
C225 a_5743_n6391# ADC15_OUT[0] 0.01fF
C226 RWLB[0] RWLB[2] 0.02fF
C227 m1_1095_5034# Din[2] 0.00fF
C228 ADC6_OUT[2] ADC7_OUT[3] 0.01fF
C229 a_5632_n6430# ADC12_OUT[1] 0.01fF
C230 WWL[2] WWL[5] 0.01fF
C231 PRE_A ADC10_OUT[0] 0.00fF
C232 PRE_CLSA ADC8_OUT[0] 0.11fF
C233 RWL[2] RWLB[4] 0.01fF
C234 RWL[3] RWLB[3] 0.08fF
C235 WWL[3] WWL[4] 0.09fF
C236 EN ADC9_OUT[0] 0.00fF
C237 RWLB[2] RWL[4] 0.02fF
C238 VDD WWL[9] 0.69fF
C239 ADC3_OUT[0] ADC4_OUT[0] 0.01fF
C240 SAEN ADC15_OUT[3] 0.01fF
C241 m1_3393_5034# VDD 0.06fF
C242 ADC13_OUT[0] VCLP 0.91fF
C243 a_5743_n6391# ADC12_OUT[2] 0.94fF
C244 ADC14_OUT[0] ADC15_OUT[0] 0.02fF
C245 WWL[4] RWLB[6] 0.01fF
C246 RWL[4] RWL[6] 0.02fF
C247 VDD RWLB[12] 2.06fF
C248 WWL[5] RWLB[5] 21.69fF
C249 RWLB[4] WWL[6] 0.02fF
C250 PRE_CLSA Iref2 0.00fF
C251 m1_5694_5034# Din[10] 0.00fF
C252 VCLP Iref1 0.15fF
C253 WWL[6] RWL[8] 0.01fF
C254 RWLB[5] RWLB[8] 0.00fF
C255 WWL[7] RWL[7] 22.38fF
C256 RWLB[6] RWLB[7] 0.09fF
C257 VDD WWLD[5] 0.73fF
C258 RWL[6] WWL[8] 0.01fF
C259 VCLP ADC10_OUT[2] 0.02fF
C260 ADC3_OUT[1] ADC4_OUT[2] 0.01fF
C261 ADC4_OUT[0] ADC5_OUT[3] 0.00fF
C262 PRE_CLSA ADC10_OUT[3] 0.10fF
C263 ADC13_OUT[0] ADC13_OUT[2] 0.03fF
C264 ADC8_OUT[1] Iref1 0.01fF
C265 SAEN ADC9_OUT[2] 0.01fF
C266 ADC10_OUT[0] Iref2 0.01fF
C267 WWL[8] WWL[10] 0.03fF
C268 RWLB[7] RWL[10] 0.01fF
C269 VDD SA_OUT[7] 1.19fF
C270 RWL[8] RWLB[9] 0.01fF
C271 RWLB[8] RWL[9] 1.23fF
C272 RWL[7] RWLB[10] 0.00fF
C273 VDD ADC8_OUT[2] 1.52fF
C274 ADC13_OUT[1] Iref2 0.01fF
C275 ADC14_OUT[1] ADC15_OUT[2] 0.01fF
C276 ADC10_OUT[0] ADC10_OUT[3] 0.03fF
C277 ADC9_OUT[1] ADC9_OUT[2] 3.83fF
C278 VDD ADC13_OUT[3] 1.58fF
C279 WWL[10] RWLB[11] 0.01fF
C280 WWL[9] RWLB[12] 0.00fF
C281 RWL[9] RWL[12] 0.00fF
C282 PRE_SRAM Din[0] 0.01fF
C283 VDD Din[1] 0.26fF
C284 RWLB[9] WWL[12] 0.00fF
C285 RWL[10] RWL[11] 0.09fF
C286 RWLB[10] WWL[11] 0.02fF
C287 m1_2243_5034# PRE_SRAM 0.14fF
C288 ADC1_OUT[2] Iref3 0.01fF
C289 Iref2 ADC1_OUT[3] 0.00fF
C290 ADC11_OUT[0] SAEN 0.06fF
C291 ADC11_OUT[2] ADC12_OUT[2] 0.01fF
C292 ADC11_OUT[1] ADC12_OUT[3] 0.00fF
C293 WWLD[3] Din[7] 0.00fF
C294 WWLD[2] Din[8] 0.00fF
C295 WWL[12] RWL[13] 0.02fF
C296 RWL[11] WWL[14] 0.00fF
C297 WWL[1] Din[3] 0.00fF
C298 RWLB[11] RWLB[13] 0.02fF
C299 RWL[12] WWL[13] 0.01fF
C300 WWLD[1] Din[9] 0.00fF
C301 RWL[0] Din[5] 0.00fF
C302 RWLB[1] Din[1] 0.01fF
C303 WWL[2] Din[0] 0.00fF
C304 PRE_SRAM Din[11] 0.01fF
C305 VDD Din[12] 0.29fF
C306 WWLD[0] Din[10] 0.00fF
C307 WWL[11] RWL[14] 0.00fF
C308 WWL[0] Din[6] 0.00fF
C309 RWLB[0] Din[4] 0.01fF
C310 RWL[1] Din[2] 0.00fF
C311 SAEN ADC14_OUT[1] 0.03fF
C312 ADC5_OUT[3] ADC6_OUT[3] 0.02fF
C313 ADC5_OUT[0] SAEN 0.07fF
C314 ADC4_OUT[0] Iref0 0.03fF
C315 ADC1_OUT[0] ADC2_OUT[1] 0.00fF
C316 PRE_CLSA ADC4_OUT[1] 0.10fF
C317 ADC6_OUT[0] VCLP 0.89fF
C318 WWL[2] Din[11] 0.00fF
C319 RWLB[13] RWL[15] 0.01fF
C320 RWL[3] Din[7] 0.00fF
C321 WWL[14] WWL[15] 0.10fF
C322 RWL[13] RWLB[15] 0.01fF
C323 RWL[5] Din[1] 0.00fF
C324 WWL[4] Din[5] 0.00fF
C325 RWLB[3] Din[6] 0.01fF
C326 WWL[3] Din[8] 0.00fF
C327 WWL[1] Din[14] 0.00fF
C328 RWLB[1] Din[12] 0.01fF
C329 VDD ADC4_OUT[0] 2.27fF
C330 RWL[2] Din[10] 0.00fF
C331 RWL[4] Din[4] 0.00fF
C332 RWLB[0] Din[15] 0.01fF
C333 WWL[5] Din[2] 0.00fF
C334 RWLB[2] Din[9] 0.01fF
C335 RWLB[5] Din[0] 0.00fF
C336 RWLB[4] Din[3] 0.01fF
C337 WWL[13] WWLD[4] 0.01fF
C338 RWL[14] RWLB[14] 0.08fF
C339 RWL[1] Din[13] 0.00fF
C340 m1_3968_5034# Din[6] 0.00fF
C341 ADC7_OUT[0] ADC7_OUT[1] 5.52fF
C342 WWL[15] SA_OUT[0] 0.08fF
C343 WWL[6] Din[10] 0.00fF
C344 RWLB[7] Din[5] 0.01fF
C345 WWL[7] Din[7] 0.00fF
C346 RWLB[5] Din[11] 0.01fF
C347 RWLB[6] Din[8] 0.01fF
C348 WWL[8] Din[4] 0.00fF
C349 RWL[8] Din[3] 0.00fF
C350 RWL[6] Din[9] 0.00fF
C351 RWLB[4] Din[14] 0.01fF
C352 RWL[4] Din[15] 0.00fF
C353 RWL[9] Din[0] 0.00fF
C354 WWL[9] Din[1] 0.00fF
C355 RWL[7] Din[6] 0.00fF
C356 RWL[5] Din[12] 0.00fF
C357 RWLB[8] Din[2] 0.01fF
C358 WWLD[4] WWLD[6] 0.03fF
C359 WWL[5] Din[13] 0.00fF
C360 a_5743_n6391# ADC7_OUT[0] 0.00fF
C361 SA_OUT[0] SA_OUT[3] 0.00fF
C362 RWL[12] Din[2] 0.00fF
C363 WWLD[5] SA_OUT[7] 0.00fF
C364 WWL[8] Din[15] 0.00fF
C365 SA_OUT[1] SA_OUT[2] 4.54fF
C366 RWLB[9] Din[10] 0.01fF
C367 WWLD[6] SA_OUT[6] 0.01fF
C368 RWLB[11] Din[4] 0.01fF
C369 WWL[11] Din[6] 0.00fF
C370 WWL[13] Din[0] 0.00fF
C371 WWL[12] Din[3] 0.00fF
C372 RWL[11] Din[5] 0.00fF
C373 WWL[10] Din[9] 0.00fF
C374 RWLB[8] Din[13] 0.01fF
C375 RWLB[10] Din[7] 0.01fF
C376 WWLD[7] SA_OUT[5] 0.05fF
C377 RWL[8] Din[14] 0.00fF
C378 RWL[10] Din[8] 0.00fF
C379 WWL[9] Din[12] 0.00fF
C380 RWL[9] Din[11] 0.00fF
C381 RWLB[12] Din[1] 0.01fF
C382 PRE_VLSA SA_OUT[4] 0.22fF
C383 ADC2_OUT[2] ADC3_OUT[2] 0.01fF
C384 VCLP ADC8_OUT[3] 1.01fF
C385 ADC2_OUT[1] ADC3_OUT[3] 0.00fF
C386 ADC6_OUT[1] Iref2 0.01fF
C387 ADC8_OUT[0] Iref3 0.01fF
C388 SAEN ADC7_OUT[3] 0.02fF
C389 m1_8567_5034# Din[14] 0.00fF
C390 VDD ADC6_OUT[3] 1.57fF
C391 Iref0 ADC12_OUT[1] 0.00fF
C392 m1_7418_5034# m1_7993_5034# 0.00fF
C393 a_5632_n6430# ADC9_OUT[2] 0.02fF
C394 WWL[12] Din[14] 0.00fF
C395 RWL[12] Din[13] 0.00fF
C396 WWL[14] Din[8] 0.00fF
C397 SA_OUT[6] SA_OUT[8] 0.03fF
C398 RWLB[12] Din[12] 0.01fF
C399 RWL[15] Din[4] 0.00fF
C400 SA_OUT[4] SA_OUT[10] 0.01fF
C401 RWLB[11] Din[15] 0.01fF
C402 WWLD[6] Din[0] 0.00fF
C403 SA_OUT[5] SA_OUT[9] 0.01fF
C404 WWLD[5] Din[1] 0.00fF
C405 SA_OUT[0] SA_OUT[14] 0.00fF
C406 RWLB[14] Din[6] 0.01fF
C407 RWL[14] Din[7] 0.00fF
C408 RWLB[13] Din[9] 0.01fF
C409 WWL[15] Din[5] 0.00fF
C410 SA_OUT[2] SA_OUT[12] 0.01fF
C411 RWLB[15] Din[3] 0.01fF
C412 WWLD[4] Din[2] 0.00fF
C413 RWL[13] Din[10] 0.00fF
C414 WWL[13] Din[11] 0.00fF
C415 PRE_VLSA SA_OUT[15] 0.11fF
C416 SA_OUT[3] SA_OUT[11] 0.01fF
C417 SA_OUT[1] SA_OUT[13] 0.00fF
C418 VDD ADC12_OUT[1] 1.57fF
C419 ADC8_OUT[1] ADC8_OUT[3] 0.01fF
C420 Iref2 Iref3 10.18fF
C421 RWL[15] Din[15] 0.00fF
C422 SA_OUT[10] SA_OUT[15] 0.02fF
C423 RWLB[15] Din[14] 0.01fF
C424 SA_OUT[1] Din[7] 0.01fF
C425 PRE_VLSA Din[9] 0.02fF
C426 SA_OUT[2] Din[6] 0.01fF
C427 SA_OUT[11] SA_OUT[14] 0.01fF
C428 SA_OUT[12] SA_OUT[13] 3.70fF
C429 SA_OUT[4] Din[4] 0.00fF
C430 WWLD[5] Din[12] 0.00fF
C431 SA_OUT[9] WE 0.02fF
C432 WWLD[6] Din[11] 0.00fF
C433 SA_OUT[3] Din[5] 0.01fF
C434 WWLD[7] Din[10] 0.00fF
C435 WWLD[4] Din[13] 0.00fF
C436 SA_OUT[0] Din[8] 0.02fF
C437 a_5632_n6430# ADC11_OUT[0] 0.01fF
C438 ADC10_OUT[3] Iref3 0.01fF
C439 SA_OUT[7] Din[12] 0.01fF
C440 SA_OUT[6] Din[13] 0.01fF
C441 SA_OUT[9] Din[10] 0.01fF
C442 SA_OUT[4] Din[15] 0.01fF
C443 SA_OUT[8] Din[11] 0.01fF
C444 WE Din[3] 0.01fF
C445 SA_OUT[5] Din[14] 0.01fF
C446 SA_OUT[3] PRE_A 0.00fF
C447 SA_OUT[2] EN 0.00fF
C448 SAEN ADC1_OUT[1] 0.04fF
C449 VCLP ADC2_OUT[1] 0.91fF
C450 ADC2_OUT[0] Iref1 0.02fF
C451 PRE_CLSA ADC2_OUT[2] 0.09fF
C452 ADC0_OUT[0] ADC1_OUT[2] 0.00fF
C453 a_5632_n6430# ADC14_OUT[1] 0.01fF
C454 VDD ADC0_OUT[1] 1.53fF
C455 SA_OUT[14] PRE_A 0.04fF
C456 SA_OUT[15] Din[15] 0.00fF
C457 Din[6] Din[7] 0.02fF
C458 VDD PRE_SRAM 6.60fF
C459 SA_OUT[13] EN 0.00fF
C460 WE Din[14] 0.01fF
C461 ADC6_OUT[0] ADC6_OUT[2] 0.03fF
C462 m1_4543_5034# VDD 0.06fF
C463 ADC15_OUT[0] VCLP 0.77fF
C464 a_5743_n6391# ADC14_OUT[2] 0.92fF
C465 WWLD[3] RWL[0] 0.94fF
C466 VDD WWL[2] 0.69fF
C467 Din[8] PRE_A 0.00fF
C468 Din[7] EN 0.02fF
C469 WWLD[2] RWLB[0] 0.01fF
C470 ADC1_OUT[2] ADC2_OUT[3] 0.01fF
C471 ADC4_OUT[1] Iref3 0.01fF
C472 ADC4_OUT[2] Iref2 0.02fF
C473 RWL[1] RWL[2] 0.09fF
C474 EN PRE_CLSA 0.04fF
C475 WWL[1] RWLB[2] 0.01fF
C476 RWL[0] RWL[3] 0.00fF
C477 RWLB[0] WWL[3] 0.01fF
C478 RWLB[1] WWL[2] 0.02fF
C479 WWL[0] RWLB[3] 0.00fF
C480 PRE_A ADC0_OUT[0] 0.00fF
C481 VDD RWLB[5] 2.06fF
C482 VCLP ADC12_OUT[2] 0.02fF
C483 PRE_CLSA ADC12_OUT[3] 0.10fF
C484 ADC14_OUT[0] ADC14_OUT[2] 0.03fF
C485 ADC12_OUT[0] Iref2 0.01fF
C486 ADC7_OUT[2] ADC7_OUT[3] 1.34fF
C487 WWL[3] RWL[4] 0.03fF
C488 Iref0 ADC15_OUT[3] 1.04fF
C489 ADC15_OUT[1] Iref2 0.01fF
C490 WWL[2] RWL[5] 0.00fF
C491 RWL[3] WWL[4] 0.01fF
C492 VDD RWL[9] 2.83fF
C493 Iref1 ADC15_OUT[2] 0.00fF
C494 EN ADC10_OUT[0] 0.00fF
C495 RWL[2] WWL[5] 0.00fF
C496 PRE_CLSA ADC9_OUT[0] 0.11fF
C497 RWLB[2] RWLB[4] 0.02fF
C498 ADC11_OUT[0] ADC11_OUT[3] 0.03fF
C499 VDD ADC15_OUT[3] 1.51fF
C500 m1_3393_5034# PRE_SRAM 0.14fF
C501 ADC13_OUT[0] SAEN 0.06fF
C502 WWL[5] WWL[6] 0.10fF
C503 VDD WWL[13] 0.69fF
C504 RWLB[4] RWL[6] 0.01fF
C505 WWL[4] WWL[7] 0.01fF
C506 ADC12_OUT[1] ADC13_OUT[3] 0.00fF
C507 ADC9_OUT[0] ADC10_OUT[0] 0.01fF
C508 ADC12_OUT[2] ADC13_OUT[2] 0.01fF
C509 RWL[5] RWLB[5] 0.08fF
C510 RWL[4] RWLB[6] 0.01fF
C511 VCLP ADC0_OUT[2] 0.95fF
C512 PRE_CLSA ADC0_OUT[3] 0.13fF
C513 SAEN Iref1 0.16fF
C514 ADC0_OUT[0] Iref2 0.01fF
C515 WWL[7] RWLB[7] 21.69fF
C516 WWL[6] RWLB[8] 0.01fF
C517 VDD WWLD[6] 0.84fF
C518 RWLB[6] WWL[8] 0.02fF
C519 RWL[6] RWL[8] 0.02fF
C520 ADC4_OUT[1] ADC4_OUT[2] 3.80fF
C521 SAEN ADC10_OUT[2] 0.01fF
C522 ADC5_OUT[0] ADC5_OUT[3] 0.03fF
C523 ADC9_OUT[1] Iref1 0.01fF
C524 VDD SA_OUT[8] 1.20fF
C525 RWL[8] WWL[10] 0.01fF
C526 RWLB[8] RWLB[9] 0.09fF
C527 WWL[9] RWL[9] 22.38fF
C528 RWLB[7] RWLB[10] 0.00fF
C529 WWL[8] RWL[10] 0.01fF
C530 VDD ADC9_OUT[2] 1.54fF
C531 ADC9_OUT[1] ADC10_OUT[2] 0.01fF
C532 PRE_SRAM Din[1] 0.01fF
C533 RWL[10] RWLB[11] 0.01fF
C534 VDD Din[2] 0.29fF
C535 RWLB[10] RWL[11] 1.23fF
C536 WWL[10] WWL[12] 0.03fF
C537 WWLD[0] Din[0] 0.00fF
C538 RWLB[9] RWL[12] 0.01fF
C539 ADC0_OUT[3] ADC1_OUT[3] 0.02fF
C540 PRE_CLSA ADC11_OUT[1] 0.10fF
C541 Iref2 ADC2_OUT[3] 0.00fF
C542 ADC11_OUT[0] Iref0 0.03fF
C543 ADC2_OUT[2] Iref3 0.01fF
C544 VDD ADC11_OUT[0] 2.27fF
C545 RWLB[1] Din[2] 0.01fF
C546 RWL[11] RWL[14] 0.00fF
C547 PRE_SRAM Din[12] 0.01fF
C548 WWL[1] Din[4] 0.00fF
C549 VDD Din[13] 0.26fF
C550 WWL[11] RWLB[14] 0.00fF
C551 WWL[2] Din[1] 0.00fF
C552 RWL[12] RWL[13] 0.09fF
C553 WWL[0] Din[7] 0.00fF
C554 RWL[2] Din[0] 0.00fF
C555 RWLB[0] Din[5] 0.01fF
C556 RWLB[11] WWL[14] 0.00fF
C557 WWL[12] RWLB[13] 0.01fF
C558 RWL[0] Din[6] 0.00fF
C559 WWLD[3] Din[8] 0.00fF
C560 RWL[1] Din[3] 0.00fF
C561 WWLD[1] Din[10] 0.00fF
C562 WWLD[2] Din[9] 0.00fF
C563 RWLB[12] WWL[13] 0.02fF
C564 WWLD[0] Din[11] 0.00fF
C565 m1_7993_5034# m1_8567_5034# 0.00fF
C566 Iref0 ADC14_OUT[1] 0.00fF
C567 ADC10_OUT[0] ADC11_OUT[1] 0.00fF
C568 ADC5_OUT[0] Iref0 0.03fF
C569 ADC6_OUT[0] SAEN 0.07fF
C570 PRE_CLSA ADC5_OUT[1] 0.10fF
C571 ADC7_OUT[0] VCLP 0.87fF
C572 ADC2_OUT[0] ADC2_OUT[1] 5.46fF
C573 VDD ADC14_OUT[1] 1.62fF
C574 RWL[5] Din[2] 0.00fF
C575 RWLB[3] Din[7] 0.01fF
C576 WWL[1] Din[15] 0.00fF
C577 RWL[1] Din[14] 0.00fF
C578 RWLB[1] Din[13] 0.01fF
C579 RWL[14] WWL[15] 0.01fF
C580 RWL[4] Din[5] 0.00fF
C581 WWL[14] RWL[15] 0.02fF
C582 WWL[3] Din[9] 0.00fF
C583 RWLB[2] Din[10] 0.01fF
C584 RWLB[5] Din[1] 0.01fF
C585 WWL[2] Din[12] 0.00fF
C586 WWL[5] Din[3] 0.00fF
C587 RWLB[13] RWLB[15] 0.02fF
C588 RWL[3] Din[8] 0.00fF
C589 WWL[4] Din[6] 0.00fF
C590 RWL[2] Din[11] 0.00fF
C591 VDD ADC5_OUT[0] 2.26fF
C592 WWL[6] Din[0] 0.00fF
C593 RWLB[4] Din[4] 0.01fF
C594 RWL[13] WWLD[4] 0.00fF
C595 m1_3968_5034# Din[7] 0.00fF
C596 ADC7_OUT[0] ADC8_OUT[1] 0.00fF
C597 RWL[7] Din[7] 0.00fF
C598 RWLB[9] Din[0] 0.00fF
C599 RWL[15] SA_OUT[0] 0.04fF
C600 RWL[5] Din[13] 0.00fF
C601 a_5632_n6430# ADC13_OUT[0] 0.01fF
C602 WWLD[5] WWLD[6] 0.69fF
C603 RWL[9] Din[1] 0.00fF
C604 WWL[6] Din[11] 0.00fF
C605 WWL[9] Din[2] 0.00fF
C606 RWLB[7] Din[6] 0.01fF
C607 RWL[8] Din[4] 0.00fF
C608 RWLB[8] Din[3] 0.01fF
C609 WWL[7] Din[8] 0.00fF
C610 RWLB[5] Din[12] 0.01fF
C611 RWLB[4] Din[15] 0.01fF
C612 RWL[6] Din[10] 0.00fF
C613 WWL[15] SA_OUT[1] 0.01fF
C614 WWL[8] Din[5] 0.00fF
C615 WWL[5] Din[14] 0.00fF
C616 RWLB[6] Din[9] 0.01fF
C617 WWLD[4] WWLD[7] 0.00fF
C618 a_5743_n6391# ADC8_OUT[0] 0.02fF
C619 ADC12_OUT[3] Iref3 0.01fF
C620 a_5632_n6430# Iref1 0.00fF
C621 WWL[13] Din[1] 0.00fF
C622 WWL[10] Din[10] 0.00fF
C623 RWL[8] Din[15] 0.00fF
C624 WWL[9] Din[13] 0.00fF
C625 RWLB[10] Din[8] 0.01fF
C626 RWL[9] Din[12] 0.00fF
C627 RWLB[9] Din[11] 0.01fF
C628 SA_OUT[0] SA_OUT[4] 0.00fF
C629 RWL[10] Din[9] 0.00fF
C630 WWLD[7] SA_OUT[6] 0.04fF
C631 RWL[13] Din[0] 0.00fF
C632 RWLB[12] Din[2] 0.01fF
C633 WWLD[6] SA_OUT[7] 0.01fF
C634 WWL[12] Din[4] 0.00fF
C635 PRE_VLSA SA_OUT[5] 0.25fF
C636 RWLB[8] Din[14] 0.01fF
C637 RWL[12] Din[3] 0.01fF
C638 SA_OUT[1] SA_OUT[3] 0.01fF
C639 RWL[11] Din[6] 0.00fF
C640 WWL[11] Din[7] 0.00fF
C641 WWLD[5] SA_OUT[8] 0.00fF
C642 RWLB[11] Din[5] 0.01fF
C643 VCLP ADC9_OUT[3] 1.03fF
C644 ADC9_OUT[0] Iref3 0.01fF
C645 ADC3_OUT[1] ADC3_OUT[3] 0.01fF
C646 ADC7_OUT[1] Iref2 0.01fF
C647 SAEN ADC8_OUT[3] 0.02fF
C648 m1_8567_5034# Din[15] 0.00fF
C649 m1_5694_5034# VDD 0.06fF
C650 VDD ADC7_OUT[3] 1.57fF
C651 a_5632_n6430# ADC10_OUT[2] 0.02fF
C652 a_5743_n6391# Iref2 0.06fF
C653 SA_OUT[5] SA_OUT[10] 0.01fF
C654 PRE_VLSA WE 2.12fF
C655 WWLD[5] Din[2] 0.00fF
C656 RWLB[14] Din[7] 0.01fF
C657 RWLB[13] Din[10] 0.01fF
C658 SA_OUT[6] SA_OUT[9] 0.03fF
C659 RWL[14] Din[8] 0.00fF
C660 RWL[12] Din[14] 0.00fF
C661 SA_OUT[4] SA_OUT[11] 0.01fF
C662 SA_OUT[0] SA_OUT[15] 0.00fF
C663 SA_OUT[3] SA_OUT[12] 0.01fF
C664 WWL[13] Din[12] 0.00fF
C665 SA_OUT[1] SA_OUT[14] 0.00fF
C666 SA_OUT[7] SA_OUT[8] 5.50fF
C667 WWLD[4] Din[3] 0.00fF
C668 WWL[12] Din[15] 0.00fF
C669 WWLD[7] Din[0] 0.00fF
C670 SA_OUT[2] SA_OUT[13] 0.01fF
C671 RWLB[12] Din[13] 0.01fF
C672 RWL[15] Din[5] 0.00fF
C673 RWLB[15] Din[4] 0.01fF
C674 WWL[14] Din[9] 0.00fF
C675 WWL[15] Din[6] 0.00fF
C676 RWL[13] Din[11] 0.00fF
C677 WWLD[6] Din[1] 0.00fF
C678 ADC8_OUT[2] ADC9_OUT[2] 0.01fF
C679 ADC8_OUT[1] ADC9_OUT[3] 0.00fF
C680 SA_OUT[4] Din[5] 0.01fF
C681 WWLD[5] Din[13] 0.00fF
C682 SA_OUT[11] SA_OUT[15] 0.01fF
C683 WWLD[6] Din[12] 0.00fF
C684 SA_OUT[10] WE 0.02fF
C685 RWLB[15] Din[15] 0.01fF
C686 SA_OUT[0] Din[9] 0.02fF
C687 ADC0_OUT[3] Iref3 0.00fF
C688 PRE_VLSA Din[10] 0.02fF
C689 SA_OUT[2] Din[7] 0.01fF
C690 SA_OUT[1] Din[8] 0.01fF
C691 SA_OUT[12] SA_OUT[14] 0.01fF
C692 WWLD[7] Din[11] 0.00fF
C693 SA_OUT[3] Din[6] 0.01fF
C694 WWLD[4] Din[14] 0.00fF
C695 VCLP ADC14_OUT[2] 0.02fF
C696 ADC15_OUT[0] ADC15_OUT[2] 0.03fF
C697 PRE_CLSA ADC14_OUT[3] 0.10fF
C698 ADC14_OUT[0] Iref2 0.01fF
C699 SA_OUT[8] Din[12] 0.01fF
C700 SA_OUT[10] Din[10] 0.00fF
C701 SA_OUT[4] PRE_A 0.00fF
C702 SA_OUT[5] Din[15] 0.01fF
C703 SA_OUT[3] EN 0.00fF
C704 SA_OUT[6] Din[14] 0.01fF
C705 SA_OUT[9] Din[11] 0.01fF
C706 WE Din[4] 0.01fF
C707 SA_OUT[7] Din[13] 0.01fF
C708 Din[1] Din[2] 0.02fF
C709 m1_2243_5034# Din[3] 0.00fF
C710 Iref0 ADC1_OUT[1] 0.00fF
C711 PRE_CLSA ADC3_OUT[2] 0.09fF
C712 ADC3_OUT[0] Iref1 0.02fF
C713 VCLP ADC3_OUT[1] 0.94fF
C714 ADC1_OUT[0] ADC1_OUT[2] 0.03fF
C715 SAEN ADC2_OUT[1] 0.04fF
C716 VDD ADC1_OUT[1] 1.57fF
C717 ADC12_OUT[0] ADC12_OUT[3] 0.03fF
C718 WE Din[15] 0.01fF
C719 VDD WWLD[0] 1.18fF
C720 ADC6_OUT[0] ADC7_OUT[2] 0.00fF
C721 ADC5_OUT[1] ADC6_OUT[1] 0.01fF
C722 SA_OUT[14] EN 0.02fF
C723 SA_OUT[15] PRE_A 0.01fF
C724 m1_4543_5034# PRE_SRAM 0.14fF
C725 ADC15_OUT[0] SAEN 0.03fF
C726 ADC13_OUT[1] ADC14_OUT[3] 0.00fF
C727 ADC13_OUT[2] ADC14_OUT[2] 0.01fF
C728 ADC11_OUT[1] Iref3 0.01fF
C729 ADC11_OUT[2] Iref2 0.02fF
C730 Din[12] Din[13] 0.02fF
C731 WWLD[2] WWL[1] 0.01fF
C732 Din[8] EN 0.00fF
C733 VDD RWL[2] 2.83fF
C734 Din[9] PRE_A 0.00fF
C735 WWLD[3] RWLB[0] 0.01fF
C736 WWL[0] RWL[0] 22.38fF
C737 m1_6843_5034# Din[11] 0.00fF
C738 ADC10_OUT[2] ADC11_OUT[3] 0.01fF
C739 ADC5_OUT[1] Iref3 0.01fF
C740 ADC5_OUT[2] Iref2 0.02fF
C741 ADC2_OUT[2] ADC2_OUT[3] 1.28fF
C742 RWLB[1] RWL[2] 1.23fF
C743 RWL[0] RWLB[3] 0.00fF
C744 EN ADC0_OUT[0] 0.00fF
C745 PRE_A ADC1_OUT[0] 0.00fF
C746 RWLB[0] RWL[3] 0.01fF
C747 WWL[1] WWL[3] 0.03fF
C748 VDD WWL[6] 0.69fF
C749 RWL[1] RWLB[2] 0.01fF
C750 SAEN ADC12_OUT[2] 0.01fF
C751 ADC7_OUT[2] ADC8_OUT[3] 0.01fF
C752 RWL[2] RWL[5] 0.00fF
C753 RWL[3] RWL[4] 0.08fF
C754 PRE_CLSA ADC10_OUT[0] 0.11fF
C755 WWL[3] RWLB[4] 0.01fF
C756 RWLB[3] WWL[4] 0.02fF
C757 WWL[2] RWLB[5] 0.00fF
C758 RWLB[2] WWL[5] 0.00fF
C759 ADC4_OUT[0] ADC5_OUT[0] 0.01fF
C760 VDD RWLB[9] 2.06fF
C761 PRE_CLSA ADC13_OUT[1] 0.10fF
C762 ADC13_OUT[0] Iref0 0.03fF
C763 WWL[5] RWL[6] 0.02fF
C764 RWLB[4] RWLB[6] 0.02fF
C765 RWL[4] WWL[7] 0.00fF
C766 WWL[4] RWL[7] 0.01fF
C767 VDD RWL[13] 2.83fF
C768 RWL[5] WWL[6] 0.01fF
C769 VDD ADC13_OUT[0] 2.28fF
C770 ADC1_OUT[0] Iref2 0.01fF
C771 ADC0_OUT[0] ADC0_OUT[3] 0.03fF
C772 m1_8567_5034# m1_9142_5034# 0.00fF
C773 VCLP ADC1_OUT[2] 0.96fF
C774 PRE_CLSA ADC1_OUT[3] 0.10fF
C775 Iref0 Iref1 13.73fF
C776 SAEN ADC0_OUT[2] 0.05fF
C777 ADC11_OUT[0] ADC12_OUT[1] 0.00fF
C778 RWL[7] RWLB[7] 0.08fF
C779 VDD WWLD[7] 1.14fF
C780 RWLB[6] RWL[8] 0.01fF
C781 WWL[6] WWL[9] 0.01fF
C782 WWL[7] WWL[8] 0.10fF
C783 RWL[6] RWLB[8] 0.01fF
C784 VDD Iref1 0.42fF
C785 ADC5_OUT[0] ADC6_OUT[3] 0.00fF
C786 ADC4_OUT[1] ADC5_OUT[2] 0.01fF
C787 ADC10_OUT[1] Iref1 0.01fF
C788 WWL[9] RWLB[9] 21.69fF
C789 RWL[8] RWL[10] 0.02fF
C790 VDD SA_OUT[9] 1.23fF
C791 RWLB[8] WWL[10] 0.02fF
C792 WWL[8] RWLB[10] 0.01fF
C793 VDD ADC10_OUT[2] 1.53fF
C794 a_5632_n6430# ADC15_OUT[0] 0.01fF
C795 ADC10_OUT[1] ADC10_OUT[2] 3.85fF
C796 WWLD[0] Din[1] 0.00fF
C797 ADC14_OUT[3] Iref3 0.01fF
C798 RWL[10] WWL[12] 0.01fF
C799 RWLB[9] RWLB[12] 0.00fF
C800 WWL[11] RWL[11] 22.38fF
C801 WWLD[1] Din[0] 0.00fF
C802 RWLB[10] RWLB[11] 0.09fF
C803 PRE_SRAM Din[2] 0.01fF
C804 WWL[10] RWL[12] 0.02fF
C805 VDD Din[3] 0.26fF
C806 Iref2 ADC3_OUT[3] 0.00fF
C807 m1_519_5034# m1_1095_5034# 0.00fF
C808 ADC3_OUT[2] Iref3 0.01fF
C809 WWL[0] Din[8] 0.00fF
C810 RWL[0] Din[7] 0.00fF
C811 RWL[2] Din[1] 0.00fF
C812 RWLB[2] Din[0] 0.00fF
C813 WWLD[2] Din[10] 0.00fF
C814 WWLD[3] Din[9] 0.00fF
C815 VDD Din[14] 0.29fF
C816 WWLD[0] Din[12] 0.00fF
C817 RWLB[11] RWL[14] 0.01fF
C818 RWLB[0] Din[6] 0.01fF
C819 RWL[12] RWLB[13] 0.01fF
C820 WWL[12] WWL[14] 0.03fF
C821 PRE_SRAM Din[13] 0.01fF
C822 RWL[1] Din[4] 0.00fF
C823 WWL[1] Din[5] 0.00fF
C824 RWLB[1] Din[3] 0.01fF
C825 WWLD[1] Din[11] 0.00fF
C826 RWLB[12] RWL[13] 1.23fF
C827 WWL[2] Din[2] 0.00fF
C828 m1_6843_5034# VDD 0.06fF
C829 ADC6_OUT[3] ADC7_OUT[3] 0.02fF
C830 a_5632_n6430# ADC12_OUT[2] 0.02fF
C831 ADC8_OUT[0] VCLP 0.86fF
C832 ADC2_OUT[0] ADC3_OUT[1] 0.00fF
C833 ADC7_OUT[0] SAEN 0.07fF
C834 ADC6_OUT[0] Iref0 0.03fF
C835 PRE_CLSA ADC6_OUT[1] 0.10fF
C836 WWL[2] Din[13] 0.00fF
C837 RWLB[5] Din[2] 0.01fF
C838 WWL[4] Din[7] 0.00fF
C839 VDD ADC6_OUT[0] 2.27fF
C840 RWLB[1] Din[14] 0.01fF
C841 RWL[2] Din[12] 0.00fF
C842 RWL[14] RWL[15] 0.09fF
C843 RWL[3] Din[9] 0.00fF
C844 RWLB[13] WWLD[4] 0.01fF
C845 RWL[4] Din[6] 0.00fF
C846 WWL[6] Din[1] 0.00fF
C847 RWLB[2] Din[11] 0.01fF
C848 RWLB[4] Din[5] 0.01fF
C849 WWL[5] Din[4] 0.00fF
C850 RWL[6] Din[0] 0.00fF
C851 RWL[1] Din[15] 0.00fF
C852 RWLB[3] Din[8] 0.01fF
C853 RWLB[14] WWL[15] 0.02fF
C854 WWL[3] Din[10] 0.00fF
C855 RWL[5] Din[3] 0.00fF
C856 WWL[14] RWLB[15] 0.01fF
C857 ADC8_OUT[0] ADC8_OUT[1] 5.52fF
C858 WWL[8] Din[6] 0.00fF
C859 RWL[5] Din[14] 0.00fF
C860 RWLB[5] Din[13] 0.01fF
C861 WWLD[5] WWLD[7] 0.03fF
C862 WWL[7] Din[9] 0.00fF
C863 WWL[5] Din[15] 0.00fF
C864 RWLB[6] Din[10] 0.01fF
C865 RWLB[8] Din[4] 0.01fF
C866 RWL[7] Din[8] 0.00fF
C867 RWLB[15] SA_OUT[0] 0.07fF
C868 RWLB[9] Din[1] 0.01fF
C869 WWL[6] Din[12] 0.00fF
C870 RWLB[7] Din[7] 0.01fF
C871 RWL[9] Din[2] 0.00fF
C872 RWL[15] SA_OUT[1] 0.00fF
C873 RWL[8] Din[5] 0.00fF
C874 RWL[6] Din[11] 0.00fF
C875 WWL[10] Din[0] 0.00fF
C876 WWL[9] Din[3] 0.00fF
C877 a_5743_n6391# ADC9_OUT[0] 0.02fF
C878 PRE_CLSA Iref3 0.00fF
C879 VCLP Iref2 0.08fF
C880 RWLB[10] Din[9] 0.01fF
C881 RWL[13] Din[1] 0.00fF
C882 RWLB[11] Din[6] 0.01fF
C883 SA_OUT[0] SA_OUT[5] 0.00fF
C884 SA_OUT[1] SA_OUT[4] 0.00fF
C885 WWL[12] Din[5] 0.00fF
C886 RWLB[8] Din[15] 0.01fF
C887 WWL[10] Din[11] 0.00fF
C888 RWL[11] Din[7] 0.00fF
C889 RWLB[12] Din[3] 0.01fF
C890 SA_OUT[2] SA_OUT[3] 5.21fF
C891 WWL[9] Din[14] 0.00fF
C892 WWLD[6] SA_OUT[8] 0.00fF
C893 WWL[11] Din[8] 0.00fF
C894 PRE_VLSA SA_OUT[6] 0.25fF
C895 WWL[13] Din[2] 0.00fF
C896 WWLD[7] SA_OUT[7] 0.03fF
C897 RWL[9] Din[13] 0.00fF
C898 RWL[12] Din[4] 0.00fF
C899 RWLB[9] Din[12] 0.01fF
C900 RWLB[13] Din[0] 0.00fF
C901 RWL[10] Din[10] 0.00fF
C902 WWLD[5] SA_OUT[9] 0.00fF
C903 ADC3_OUT[1] ADC4_OUT[3] 0.00fF
C904 VCLP ADC10_OUT[3] 1.02fF
C905 SAEN ADC9_OUT[3] 0.02fF
C906 ADC10_OUT[0] Iref3 0.01fF
C907 ADC3_OUT[2] ADC4_OUT[2] 0.01fF
C908 ADC13_OUT[0] ADC13_OUT[3] 0.03fF
C909 ADC8_OUT[1] Iref2 0.01fF
C910 m1_5694_5034# PRE_SRAM 0.14fF
C911 VDD ADC8_OUT[3] 1.57fF
C912 SA_OUT[5] SA_OUT[11] 0.01fF
C913 SA_OUT[1] SA_OUT[15] 0.00fF
C914 WWLD[7] Din[1] 0.00fF
C915 SA_OUT[3] SA_OUT[13] 0.01fF
C916 RWLB[13] Din[11] 0.01fF
C917 ADC14_OUT[1] ADC15_OUT[3] 0.00fF
C918 RWLB[15] Din[5] 0.01fF
C919 WWL[15] Din[7] 0.00fF
C920 WWL[14] Din[10] 0.00fF
C921 RWL[13] Din[12] 0.00fF
C922 ADC13_OUT[1] Iref3 0.01fF
C923 SA_OUT[7] SA_OUT[9] 0.02fF
C924 SA_OUT[0] WE 0.01fF
C925 WWLD[4] Din[4] 0.00fF
C926 PRE_VLSA Din[0] 0.02fF
C927 WWLD[6] Din[2] 0.00fF
C928 ADC13_OUT[2] Iref2 0.02fF
C929 SA_OUT[4] SA_OUT[12] 0.01fF
C930 RWLB[14] Din[8] 0.01fF
C931 RWL[12] Din[15] 0.00fF
C932 ADC14_OUT[2] ADC15_OUT[2] 0.02fF
C933 WWL[13] Din[13] 0.00fF
C934 RWLB[12] Din[14] 0.01fF
C935 SA_OUT[6] SA_OUT[10] 0.03fF
C936 WWLD[5] Din[3] 0.00fF
C937 ADC15_OUT[1] ADC14_OUT[3] 0.00fF
C938 RWL[14] Din[9] 0.00fF
C939 SA_OUT[2] SA_OUT[14] 0.01fF
C940 RWL[15] Din[6] 0.00fF
C941 ADC9_OUT[1] ADC9_OUT[3] 0.01fF
C942 ADC1_OUT[3] Iref3 0.01fF
C943 SA_OUT[0] Din[10] 0.02fF
C944 WWLD[5] Din[14] 0.00fF
C945 SA_OUT[4] Din[6] 0.01fF
C946 SA_OUT[11] WE 0.02fF
C947 WWLD[7] Din[12] 0.00fF
C948 SA_OUT[2] Din[8] 0.01fF
C949 SA_OUT[3] Din[7] 0.01fF
C950 WWLD[4] Din[15] 0.00fF
C951 SA_OUT[1] Din[9] 0.01fF
C952 SA_OUT[12] SA_OUT[15] 0.01fF
C953 SA_OUT[13] SA_OUT[14] 1.17fF
C954 WWLD[6] Din[13] 0.00fF
C955 ADC11_OUT[2] ADC12_OUT[3] 0.01fF
C956 SA_OUT[5] Din[5] 0.00fF
C957 PRE_VLSA Din[11] 0.02fF
C958 SAEN ADC14_OUT[2] 0.01fF
C959 SA_OUT[9] Din[12] 0.01fF
C960 WE Din[5] 0.01fF
C961 SA_OUT[10] Din[11] 0.01fF
C962 SA_OUT[8] Din[13] 0.01fF
C963 SA_OUT[4] EN 0.00fF
C964 SA_OUT[7] Din[14] 0.01fF
C965 SA_OUT[5] PRE_A 0.00fF
C966 SA_OUT[6] Din[15] 0.01fF
C967 ADC4_OUT[0] Iref1 0.02fF
C968 Iref0 ADC2_OUT[1] 0.00fF
C969 PRE_CLSA ADC4_OUT[2] 0.09fF
C970 m1_2243_5034# Din[4] 0.00fF
C971 ADC1_OUT[0] ADC2_OUT[2] 0.00fF
C972 VCLP ADC4_OUT[1] 0.94fF
C973 ADC0_OUT[1] ADC1_OUT[1] 0.01fF
C974 SAEN ADC3_OUT[1] 0.04fF
C975 PRE_CLSA ADC12_OUT[0] 0.11fF
C976 a_5743_n6391# ADC11_OUT[1] 0.01fF
C977 VDD ADC2_OUT[1] 1.57fF
C978 a_5632_n6430# ADC7_OUT[0] 0.01fF
C979 WE PRE_A 0.05fF
C980 Din[7] Din[8] 0.02fF
C981 VDD WWLD[1] 1.01fF
C982 PRE_SRAM WWLD[0] 0.79fF
C983 ADC7_OUT[0] ADC7_OUT[2] 0.04fF
C984 ADC15_OUT[0] Iref0 0.27fF
C985 PRE_CLSA ADC15_OUT[1] 0.07fF
C986 VDD ADC15_OUT[0] 2.29fF
C987 Din[9] EN 0.02fF
C988 VDD RWLB[2] 2.06fF
C989 WWLD[2] RWL[1] 0.01fF
C990 WWLD[3] WWL[1] 0.03fF
C991 WWL[0] RWLB[0] 21.69fF
C992 Din[10] PRE_A 0.00fF
C993 m1_6843_5034# Din[12] 0.00fF
C994 ADC12_OUT[0] ADC13_OUT[1] 0.00fF
C995 ADC6_OUT[1] Iref3 0.01fF
C996 ADC2_OUT[2] ADC3_OUT[3] 0.01fF
C997 ADC6_OUT[2] Iref2 0.02fF
C998 EN ADC1_OUT[0] 0.00fF
C999 WWL[2] RWL[2] 22.38fF
C1000 RWL[1] WWL[3] 0.01fF
C1001 RWLB[0] RWLB[3] 0.00fF
C1002 VDD RWL[6] 2.83fF
C1003 WWL[1] RWL[3] 0.01fF
C1004 PRE_CLSA ADC0_OUT[0] 0.12fF
C1005 RWLB[1] RWLB[2] 0.09fF
C1006 PRE_A ADC2_OUT[0] 0.00fF
C1007 ADC12_OUT[1] Iref1 0.01fF
C1008 VDD ADC12_OUT[2] 1.54fF
C1009 ADC8_OUT[2] ADC8_OUT[3] 1.33fF
C1010 WWL[3] WWL[5] 0.03fF
C1011 RWLB[3] RWL[4] 0.97fF
C1012 RWL[3] RWLB[4] 0.01fF
C1013 RWLB[2] RWL[5] 0.01fF
C1014 VDD WWL[10] 0.70fF
C1015 ADC11_OUT[1] ADC11_OUT[2] 3.86fF
C1016 m1_519_5034# Din[0] 0.00fF
C1017 m1_1095_5034# m1_1670_5034# 0.00fF
C1018 WWL[4] RWLB[7] 0.00fF
C1019 RWL[4] RWL[7] 0.00fF
C1020 RWL[5] RWL[6] 0.09fF
C1021 RWLB[4] WWL[7] 0.01fF
C1022 WWL[5] RWLB[6] 0.01fF
C1023 RWLB[5] WWL[6] 0.02fF
C1024 VDD RWLB[13] 2.06fF
C1025 PRE_CLSA ADC2_OUT[3] 0.10fF
C1026 ADC0_OUT[1] Iref1 0.00fF
C1027 VCLP ADC2_OUT[2] 0.95fF
C1028 m1_7993_5034# VDD 0.06fF
C1029 ADC2_OUT[0] Iref2 0.01fF
C1030 ADC0_OUT[0] ADC1_OUT[3] 0.00fF
C1031 SAEN ADC1_OUT[2] 0.04fF
C1032 a_5632_n6430# ADC14_OUT[2] 0.02fF
C1033 WWL[6] RWL[9] 0.01fF
C1034 VDD ADC0_OUT[2] 1.51fF
C1035 VDD PRE_VLSA 3.62fF
C1036 RWL[6] WWL[9] 0.00fF
C1037 RWLB[6] RWLB[8] 0.02fF
C1038 RWL[7] WWL[8] 0.01fF
C1039 WWL[7] RWL[8] 0.02fF
C1040 ADC5_OUT[1] ADC5_OUT[2] 3.82fF
C1041 ADC6_OUT[0] ADC6_OUT[3] 0.03fF
C1042 m1_5118_5034# Din[8] 0.00fF
C1043 RWLB[8] RWL[10] 0.01fF
C1044 RWL[8] RWLB[10] 0.01fF
C1045 RWL[9] RWLB[9] 0.08fF
C1046 WWL[8] WWL[11] 0.01fF
C1047 VDD SA_OUT[10] 1.25fF
C1048 WWL[9] WWL[10] 0.10fF
C1049 VDD Din[4] 0.29fF
C1050 WWLD[2] Din[0] 0.00fF
C1051 WWLD[1] Din[1] 0.00fF
C1052 WWL[10] RWLB[12] 0.01fF
C1053 PRE_SRAM Din[3] 0.01fF
C1054 RWL[10] RWL[12] 0.02fF
C1055 WWL[11] RWLB[11] 21.69fF
C1056 WWLD[0] Din[2] 0.00fF
C1057 RWLB[10] WWL[12] 0.02fF
C1058 ADC4_OUT[2] Iref3 0.01fF
C1059 Iref2 ADC4_OUT[3] 0.00fF
C1060 ADC1_OUT[3] ADC2_OUT[3] 0.02fF
C1061 VCLP ADC12_OUT[3] 1.07fF
C1062 ADC14_OUT[0] ADC14_OUT[3] 0.03fF
C1063 ADC12_OUT[0] Iref3 0.01fF
C1064 WWL[13] RWL[13] 22.38fF
C1065 WWL[1] Din[6] 0.00fF
C1066 RWLB[0] Din[7] 0.01fF
C1067 RWLB[12] RWLB[13] 0.09fF
C1068 RWL[1] Din[5] 0.00fF
C1069 WWLD[1] Din[12] 0.00fF
C1070 WWLD[2] Din[11] 0.00fF
C1071 WWL[3] Din[0] 0.00fF
C1072 RWL[0] Din[8] 0.00fF
C1073 WWL[0] Din[9] 0.00fF
C1074 WWL[2] Din[3] 0.00fF
C1075 RWL[2] Din[2] 0.00fF
C1076 RWLB[2] Din[1] 0.01fF
C1077 WWL[12] RWL[14] 0.01fF
C1078 WWLD[3] Din[10] 0.00fF
C1079 PRE_SRAM Din[14] 0.01fF
C1080 VDD Din[15] 0.27fF
C1081 RWLB[1] Din[4] 0.01fF
C1082 WWLD[0] Din[13] 0.00fF
C1083 RWL[12] WWL[14] 0.01fF
C1084 RWLB[11] RWLB[14] 0.00fF
C1085 m1_6843_5034# PRE_SRAM 0.14fF
C1086 ADC3_OUT[0] ADC3_OUT[1] 5.45fF
C1087 Iref1 ADC15_OUT[3] 0.00fF
C1088 PRE_CLSA ADC7_OUT[1] 0.10fF
C1089 ADC15_OUT[1] Iref3 0.01fF
C1090 ADC7_OUT[0] Iref0 0.03fF
C1091 ADC8_OUT[0] SAEN 0.06fF
C1092 ADC9_OUT[0] VCLP 0.89fF
C1093 ADC15_OUT[2] Iref2 0.02fF
C1094 WWL[6] Din[2] 0.00fF
C1095 WWL[5] Din[5] 0.00fF
C1096 WWL[2] Din[14] 0.00fF
C1097 RWL[6] Din[1] 0.00fF
C1098 RWLB[6] Din[0] 0.00fF
C1099 RWLB[3] Din[9] 0.01fF
C1100 WWL[14] WWLD[4] 0.03fF
C1101 RWLB[4] Din[6] 0.01fF
C1102 RWLB[1] Din[15] 0.01fF
C1103 WWL[4] Din[8] 0.00fF
C1104 RWLB[14] RWL[15] 1.23fF
C1105 RWL[2] Din[13] 0.00fF
C1106 RWL[3] Din[10] 0.00fF
C1107 RWL[5] Din[4] 0.00fF
C1108 RWL[14] RWLB[15] 0.01fF
C1109 RWL[4] Din[7] 0.01fF
C1110 RWLB[5] Din[3] 0.01fF
C1111 WWL[3] Din[11] 0.00fF
C1112 VDD ADC7_OUT[0] 2.27fF
C1113 RWLB[2] Din[12] 0.01fF
C1114 a_5743_n6391# PRE_CLSA 0.43fF
C1115 ADC12_OUT[2] ADC13_OUT[3] 0.01fF
C1116 ADC8_OUT[0] ADC9_OUT[1] 0.00fF
C1117 RWLB[8] Din[5] 0.01fF
C1118 WWL[9] Din[4] 0.00fF
C1119 RWL[8] Din[6] 0.00fF
C1120 WWL[6] Din[13] 0.00fF
C1121 RWL[7] Din[9] 0.00fF
C1122 RWLB[7] Din[8] 0.01fF
C1123 RWLB[5] Din[14] 0.01fF
C1124 RWLB[9] Din[2] 0.01fF
C1125 WWLD[5] PRE_VLSA 0.00fF
C1126 WWLD[4] SA_OUT[0] 0.16fF
C1127 RWL[6] Din[12] 0.00fF
C1128 RWLB[15] SA_OUT[1] 0.01fF
C1129 WWL[8] Din[7] 0.00fF
C1130 WWL[10] Din[1] 0.00fF
C1131 RWL[9] Din[3] 0.00fF
C1132 RWLB[6] Din[11] 0.01fF
C1133 RWL[5] Din[15] 0.00fF
C1134 RWL[10] Din[0] 0.00fF
C1135 WWL[7] Din[10] 0.00fF
C1136 WWLD[6] WWLD[7] 0.86fF
C1137 VCLP ADC0_OUT[3] 1.00fF
C1138 ADC0_OUT[0] Iref3 0.01fF
C1139 SAEN Iref2 0.08fF
C1140 a_5743_n6391# ADC10_OUT[0] 0.02fF
C1141 RWL[9] Din[14] 0.00fF
C1142 SA_OUT[0] SA_OUT[6] 0.00fF
C1143 RWL[10] Din[11] 0.00fF
C1144 WWL[14] Din[0] 0.00fF
C1145 WWL[11] Din[9] 0.00fF
C1146 PRE_CLSA ADC14_OUT[0] 0.11fF
C1147 RWLB[9] Din[13] 0.01fF
C1148 WWL[12] Din[6] 0.00fF
C1149 RWL[12] Din[5] 0.00fF
C1150 RWLB[12] Din[4] 0.01fF
C1151 RWLB[10] Din[10] 0.01fF
C1152 WWL[13] Din[3] 0.00fF
C1153 WWLD[6] SA_OUT[9] 0.00fF
C1154 RWLB[13] Din[1] 0.01fF
C1155 a_5743_n6391# ADC13_OUT[1] 0.01fF
C1156 WWLD[5] SA_OUT[10] 0.00fF
C1157 RWLB[11] Din[7] 0.01fF
C1158 WWLD[7] SA_OUT[8] 0.02fF
C1159 SA_OUT[2] SA_OUT[4] 0.01fF
C1160 WWL[10] Din[12] 0.00fF
C1161 RWL[13] Din[2] 0.00fF
C1162 PRE_VLSA SA_OUT[7] 0.31fF
C1163 WWL[9] Din[15] 0.00fF
C1164 RWL[11] Din[8] 0.00fF
C1165 SA_OUT[1] SA_OUT[5] 0.00fF
C1166 ADC9_OUT[1] Iref2 0.01fF
C1167 ADC4_OUT[1] ADC4_OUT[3] 0.01fF
C1168 SAEN ADC10_OUT[3] 0.02fF
C1169 VDD ADC9_OUT[3] 1.58fF
C1170 m1_519_5034# VDD 0.06fF
C1171 SA_OUT[0] Din[0] 0.00fF
C1172 SA_OUT[7] SA_OUT[10] 0.02fF
C1173 WWLD[4] Din[5] 0.00fF
C1174 PRE_VLSA Din[1] 0.02fF
C1175 SA_OUT[1] WE 0.01fF
C1176 RWLB[12] Din[15] 0.01fF
C1177 SA_OUT[8] SA_OUT[9] 5.40fF
C1178 WWLD[6] Din[3] 0.00fF
C1179 RWLB[14] Din[9] 0.01fF
C1180 RWL[14] Din[10] 0.00fF
C1181 SA_OUT[5] SA_OUT[12] 0.01fF
C1182 RWL[15] Din[7] 0.00fF
C1183 WWL[14] Din[11] 0.00fF
C1184 SA_OUT[3] SA_OUT[14] 0.01fF
C1185 SA_OUT[4] SA_OUT[13] 0.01fF
C1186 RWLB[15] Din[6] 0.01fF
C1187 SA_OUT[2] SA_OUT[15] 0.01fF
C1188 RWLB[13] Din[12] 0.01fF
C1189 WWLD[7] Din[2] 0.00fF
C1190 SA_OUT[6] SA_OUT[11] 0.03fF
C1191 RWL[13] Din[13] 0.00fF
C1192 WWLD[5] Din[4] 0.00fF
C1193 WWL[13] Din[14] 0.00fF
C1194 WWL[15] Din[8] 0.00fF
C1195 ADC9_OUT[2] ADC10_OUT[2] 0.01fF
C1196 ADC9_OUT[1] ADC10_OUT[3] 0.00fF
C1197 SA_OUT[1] Din[10] 0.01fF
C1198 ADC13_OUT[0] ADC14_OUT[1] 0.00fF
C1199 SA_OUT[5] Din[6] 0.01fF
C1200 SA_OUT[2] Din[9] 0.01fF
C1201 VCLP ADC11_OUT[1] 0.91fF
C1202 PRE_CLSA ADC11_OUT[2] 0.09fF
C1203 SA_OUT[0] Din[11] 0.02fF
C1204 ADC2_OUT[3] Iref3 0.01fF
C1205 PRE_VLSA Din[12] 0.02fF
C1206 SA_OUT[13] SA_OUT[15] 0.01fF
C1207 ADC11_OUT[0] Iref1 0.02fF
C1208 SA_OUT[12] WE 0.02fF
C1209 WWLD[5] Din[15] 0.00fF
C1210 SA_OUT[4] Din[7] 0.01fF
C1211 WWLD[6] Din[14] 0.00fF
C1212 WWLD[7] Din[13] 0.00fF
C1213 SA_OUT[3] Din[8] 0.01fF
C1214 ADC14_OUT[1] Iref1 0.01fF
C1215 ADC10_OUT[0] ADC11_OUT[2] 0.00fF
C1216 SAEN ADC4_OUT[1] 0.04fF
C1217 PRE_CLSA ADC5_OUT[2] 0.09fF
C1218 ADC5_OUT[0] Iref1 0.02fF
C1219 Iref0 ADC3_OUT[1] 0.00fF
C1220 SA_OUT[11] Din[11] 0.00fF
C1221 SA_OUT[7] Din[15] 0.01fF
C1222 Din[2] Din[3] 0.02fF
C1223 WE Din[6] 0.01fF
C1224 VCLP ADC5_OUT[1] 0.93fF
C1225 SA_OUT[5] EN 0.00fF
C1226 SA_OUT[9] Din[13] 0.01fF
C1227 SA_OUT[8] Din[14] 0.01fF
C1228 SA_OUT[10] Din[12] 0.01fF
C1229 SA_OUT[6] PRE_A 0.00fF
C1230 ADC2_OUT[0] ADC2_OUT[2] 0.03fF
C1231 VDD ADC14_OUT[2] 1.57fF
C1232 VDD ADC3_OUT[1] 1.58fF
C1233 ADC12_OUT[1] ADC12_OUT[2] 3.83fF
C1234 a_5632_n6430# ADC8_OUT[0] 0.01fF
C1235 VDD WWLD[2] 0.74fF
C1236 Din[0] PRE_A 0.00fF
C1237 WE EN 0.10fF
C1238 PRE_SRAM WWLD[1] 0.05fF
C1239 ADC6_OUT[1] ADC7_OUT[1] 0.01fF
C1240 ADC7_OUT[0] ADC8_OUT[2] 0.00fF
C1241 m1_1670_5034# m1_2243_5034# 0.00fF
C1242 Din[11] PRE_A 0.00fF
C1243 WWL[0] WWL[1] 0.10fF
C1244 WWLD[3] RWL[1] 0.01fF
C1245 RWL[0] RWLB[0] 0.08fF
C1246 VDD WWL[3] 0.70fF
C1247 Din[10] EN 0.00fF
C1248 Din[13] Din[14] 0.02fF
C1249 WWLD[2] RWLB[1] 0.00fF
C1250 m1_9142_5034# VDD 0.06fF
C1251 a_5632_n6430# Iref2 0.08fF
C1252 ADC3_OUT[2] ADC3_OUT[3] 1.27fF
C1253 ADC7_OUT[1] Iref3 0.01fF
C1254 ADC7_OUT[2] Iref2 0.03fF
C1255 VDD RWLB[6] 2.06fF
C1256 RWL[1] RWL[3] 0.02fF
C1257 RWLB[1] WWL[3] 0.02fF
C1258 PRE_CLSA ADC1_OUT[0] 0.11fF
C1259 EN ADC2_OUT[0] 0.00fF
C1260 WWL[1] RWLB[3] 0.01fF
C1261 WWL[2] RWLB[2] 21.69fF
C1262 PRE_A ADC3_OUT[0] 0.00fF
C1263 a_5743_n6391# Iref3 0.02fF
C1264 ADC8_OUT[2] ADC9_OUT[3] 0.01fF
C1265 RWLB[2] RWLB[5] 0.00fF
C1266 RWL[3] WWL[5] 0.01fF
C1267 ADC5_OUT[0] ADC6_OUT[0] 0.01fF
C1268 WWL[4] RWL[4] 22.38fF
C1269 WWL[3] RWL[5] 0.01fF
C1270 RWLB[3] RWLB[4] 0.08fF
C1271 VDD RWL[10] 2.83fF
C1272 m1_519_5034# Din[1] 0.00fF
C1273 RWL[5] RWLB[6] 0.01fF
C1274 VDD WWL[14] 0.69fF
C1275 WWL[5] WWL[7] 0.03fF
C1276 RWLB[4] RWL[7] 0.01fF
C1277 RWLB[5] RWL[6] 1.23fF
C1278 RWL[4] RWLB[7] 0.00fF
C1279 ADC15_OUT[0] ADC15_OUT[3] 0.03fF
C1280 VCLP ADC14_OUT[3] 1.01fF
C1281 ADC14_OUT[0] Iref3 0.01fF
C1282 m1_7993_5034# PRE_SRAM 0.14fF
C1283 ADC1_OUT[1] Iref1 0.01fF
C1284 VCLP ADC3_OUT[2] 0.94fF
C1285 ADC1_OUT[0] ADC1_OUT[3] 0.03fF
C1286 PRE_CLSA ADC3_OUT[3] 0.10fF
C1287 ADC0_OUT[1] ADC0_OUT[2] 4.12fF
C1288 ADC3_OUT[0] Iref2 0.01fF
C1289 SAEN ADC2_OUT[2] 0.04fF
C1290 WWL[7] RWLB[8] 0.01fF
C1291 RWL[6] RWL[9] 0.00fF
C1292 RWLB[6] WWL[9] 0.01fF
C1293 RWLB[7] WWL[8] 0.02fF
C1294 RWL[7] RWL[8] 0.09fF
C1295 WWL[6] RWLB[9] 0.00fF
C1296 VDD SA_OUT[0] 2.69fF
C1297 VDD ADC1_OUT[2] 1.53fF
C1298 ADC5_OUT[1] ADC6_OUT[2] 0.01fF
C1299 ADC6_OUT[0] ADC7_OUT[3] 0.00fF
C1300 m1_5118_5034# Din[9] 0.00fF
C1301 WWL[8] RWL[11] 0.01fF
C1302 RWL[9] WWL[10] 0.01fF
C1303 RWLB[8] RWLB[10] 0.02fF
C1304 WWL[9] RWL[10] 0.02fF
C1305 VDD SA_OUT[11] 1.28fF
C1306 RWL[8] WWL[11] 0.00fF
C1307 ADC13_OUT[2] ADC14_OUT[3] 0.01fF
C1308 ADC11_OUT[2] Iref3 0.01fF
C1309 Iref2 ADC11_OUT[3] 0.00fF
C1310 a_5743_n6391# ADC12_OUT[0] 0.02fF
C1311 RWLB[10] RWL[12] 0.02fF
C1312 RWL[10] RWLB[12] 0.01fF
C1313 WWL[11] WWL[12] 0.09fF
C1314 ADC10_OUT[3] ADC11_OUT[3] 0.02fF
C1315 RWL[11] RWLB[11] 0.08fF
C1316 WWL[10] WWL[13] 0.01fF
C1317 PRE_SRAM Din[4] 0.01fF
C1318 VDD Din[5] 0.26fF
C1319 WWLD[3] Din[0] 0.00fF
C1320 WWLD[0] Din[3] 0.00fF
C1321 WWLD[2] Din[1] 0.00fF
C1322 WWLD[1] Din[2] 0.00fF
C1323 Iref2 ADC5_OUT[3] 0.00fF
C1324 ADC5_OUT[2] Iref3 0.01fF
C1325 a_5743_n6391# ADC15_OUT[1] 0.00fF
C1326 PRE_CLSA VCLP 7.13fF
C1327 SAEN ADC12_OUT[3] 0.02fF
C1328 RWL[12] RWL[14] 0.02fF
C1329 WWLD[0] Din[14] 0.00fF
C1330 WWL[0] Din[10] 0.00fF
C1331 WWL[3] Din[1] 0.00fF
C1332 WWL[12] RWLB[14] 0.01fF
C1333 RWL[0] Din[9] 0.00fF
C1334 PRE_SRAM Din[15] 0.01fF
C1335 WWL[13] RWLB[13] 21.69fF
C1336 RWLB[2] Din[2] 0.01fF
C1337 RWLB[1] Din[5] 0.01fF
C1338 RWL[2] Din[3] 0.00fF
C1339 WWL[1] Din[7] 0.00fF
C1340 RWLB[12] WWL[14] 0.02fF
C1341 RWL[1] Din[6] 0.00fF
C1342 VDD PRE_A 3.56fF
C1343 RWL[3] Din[0] 0.00fF
C1344 RWLB[0] Din[8] 0.01fF
C1345 WWL[2] Din[4] 0.00fF
C1346 WWLD[1] Din[13] 0.00fF
C1347 WWLD[2] Din[12] 0.00fF
C1348 WWLD[3] Din[11] 0.00fF
C1349 ADC7_OUT[3] ADC8_OUT[3] 0.02fF
C1350 m1_1670_5034# VDD 0.06fF
C1351 ADC3_OUT[0] ADC4_OUT[1] 0.00fF
C1352 ADC10_OUT[0] VCLP 0.88fF
C1353 ADC9_OUT[0] SAEN 0.06fF
C1354 PRE_CLSA ADC8_OUT[1] 0.10fF
C1355 ADC8_OUT[0] Iref0 0.03fF
C1356 RWL[3] Din[11] 0.00fF
C1357 RWLB[5] Din[4] 0.01fF
C1358 WWL[15] RWL[15] 22.38fF
C1359 RWLB[4] Din[7] 0.01fF
C1360 VDD ADC8_OUT[0] 2.27fF
C1361 WWL[5] Din[6] 0.00fF
C1362 RWLB[14] RWLB[15] 0.09fF
C1363 RWL[5] Din[5] 0.00fF
C1364 WWL[3] Din[12] 0.00fF
C1365 WWL[4] Din[9] 0.00fF
C1366 RWLB[2] Din[13] 0.01fF
C1367 RWL[4] Din[8] 0.00fF
C1368 WWL[2] Din[15] 0.00fF
C1369 RWL[14] WWLD[4] 0.01fF
C1370 WWL[7] Din[0] 0.00fF
C1371 RWLB[3] Din[10] 0.01fF
C1372 RWLB[6] Din[1] 0.01fF
C1373 RWL[6] Din[2] 0.00fF
C1374 WWL[6] Din[3] 0.00fF
C1375 RWL[2] Din[14] 0.00fF
C1376 WWL[14] WWLD[5] 0.01fF
C1377 PRE_CLSA ADC13_OUT[2] 0.09fF
C1378 ADC14_OUT[0] ADC15_OUT[1] 0.01fF
C1379 VCLP ADC13_OUT[1] 0.98fF
C1380 ADC13_OUT[0] Iref1 0.02fF
C1381 ADC9_OUT[0] ADC9_OUT[1] 5.50fF
C1382 WWL[7] Din[11] 0.00fF
C1383 RWLB[7] Din[9] 0.01fF
C1384 RWLB[6] Din[12] 0.01fF
C1385 WWL[8] Din[8] 0.00fF
C1386 RWLB[9] Din[3] 0.01fF
C1387 RWLB[8] Din[6] 0.01fF
C1388 WWLD[4] SA_OUT[1] 0.03fF
C1389 WWL[10] Din[2] 0.00fF
C1390 RWLB[10] Din[0] 0.00fF
C1391 WWL[6] Din[14] 0.00fF
C1392 RWL[10] Din[1] 0.00fF
C1393 WWL[9] Din[5] 0.00fF
C1394 RWL[8] Din[7] 0.00fF
C1395 RWL[9] Din[4] 0.00fF
C1396 WWLD[5] SA_OUT[0] 0.21fF
C1397 RWL[7] Din[10] 0.00fF
C1398 RWLB[5] Din[15] 0.01fF
C1399 WWLD[6] PRE_VLSA 0.01fF
C1400 RWL[6] Din[13] 0.00fF
C1401 VCLP ADC1_OUT[3] 1.03fF
C1402 SAEN ADC0_OUT[3] 0.02fF
C1403 Iref0 Iref2 0.01fF
C1404 ADC1_OUT[0] Iref3 0.01fF
C1405 ADC11_OUT[0] ADC12_OUT[2] 0.00fF
C1406 m1_3393_5034# Din[5] 0.00fF
C1407 VDD Iref2 0.41fF
C1408 RWLB[12] Din[5] 0.01fF
C1409 WWLD[6] SA_OUT[10] 0.00fF
C1410 RWL[14] Din[0] 0.00fF
C1411 RWLB[13] Din[2] 0.01fF
C1412 RWLB[11] Din[8] 0.01fF
C1413 SA_OUT[0] SA_OUT[7] 0.00fF
C1414 WWL[10] Din[13] 0.00fF
C1415 SA_OUT[3] SA_OUT[4] 4.44fF
C1416 RWL[9] Din[15] 0.00fF
C1417 RWLB[9] Din[14] 0.01fF
C1418 SA_OUT[2] SA_OUT[5] 0.01fF
C1419 WWL[13] Din[4] 0.00fF
C1420 RWL[13] Din[3] 0.00fF
C1421 RWL[10] Din[12] 0.00fF
C1422 RWL[11] Din[9] 0.00fF
C1423 RWLB[10] Din[11] 0.01fF
C1424 RWL[12] Din[6] 0.00fF
C1425 WWLD[5] SA_OUT[11] 0.00fF
C1426 WWLD[7] SA_OUT[9] 0.02fF
C1427 PRE_VLSA SA_OUT[8] 0.29fF
C1428 WWL[11] Din[10] 0.00fF
C1429 WWL[14] Din[1] 0.00fF
C1430 SA_OUT[1] SA_OUT[6] 0.00fF
C1431 WWL[12] Din[7] 0.00fF
C1432 ADC13_OUT[1] ADC13_OUT[2] 3.83fF
C1433 ADC10_OUT[1] Iref2 0.01fF
C1434 ADC4_OUT[2] ADC5_OUT[2] 0.01fF
C1435 ADC4_OUT[1] ADC5_OUT[3] 0.00fF
C1436 VDD ADC10_OUT[3] 1.58fF
C1437 m1_519_5034# PRE_SRAM 0.14fF
C1438 WWL[14] Din[12] 0.00fF
C1439 RWL[13] Din[14] 0.00fF
C1440 RWLB[15] Din[7] 0.01fF
C1441 RWL[15] Din[8] 0.00fF
C1442 SA_OUT[7] SA_OUT[11] 0.02fF
C1443 SA_OUT[3] SA_OUT[15] 0.01fF
C1444 RWLB[13] Din[13] 0.01fF
C1445 SA_OUT[6] SA_OUT[12] 0.03fF
C1446 SA_OUT[5] SA_OUT[13] 0.01fF
C1447 WWLD[4] Din[6] 0.00fF
C1448 WWL[13] Din[15] 0.00fF
C1449 WWLD[5] Din[5] 0.00fF
C1450 WWLD[6] Din[4] 0.00fF
C1451 RWL[14] Din[11] 0.00fF
C1452 WWLD[7] Din[3] 0.00fF
C1453 SA_OUT[0] Din[1] 0.02fF
C1454 WWL[15] Din[9] 0.00fF
C1455 m1_2243_5034# m1_2819_5034# 0.00fF
C1456 SA_OUT[2] WE 0.01fF
C1457 PRE_VLSA Din[2] 0.02fF
C1458 RWLB[14] Din[10] 0.01fF
C1459 SA_OUT[4] SA_OUT[14] 0.01fF
C1460 SA_OUT[8] SA_OUT[10] 0.02fF
C1461 ADC10_OUT[1] ADC10_OUT[3] 0.01fF
C1462 m1_7993_5034# Din[13] 0.00fF
C1463 SAEN ADC11_OUT[1] 0.03fF
C1464 WWLD[7] Din[14] 0.00fF
C1465 SA_OUT[1] Din[11] 0.01fF
C1466 WWLD[6] Din[15] 0.00fF
C1467 SA_OUT[4] Din[8] 0.01fF
C1468 SA_OUT[5] Din[7] 0.01fF
C1469 SA_OUT[2] Din[10] 0.01fF
C1470 SA_OUT[13] WE 0.10fF
C1471 SA_OUT[3] Din[9] 0.01fF
C1472 SA_OUT[14] SA_OUT[15] 1.11fF
C1473 SA_OUT[0] Din[12] 0.02fF
C1474 ADC3_OUT[3] Iref3 0.01fF
C1475 SA_OUT[6] Din[6] 0.00fF
C1476 PRE_VLSA Din[13] 0.02fF
C1477 SA_OUT[8] Din[15] 0.01fF
C1478 SA_OUT[10] Din[13] 0.01fF
C1479 SA_OUT[6] EN 0.00fF
C1480 SA_OUT[9] Din[14] 0.01fF
C1481 SA_OUT[11] Din[12] 0.01fF
C1482 WE Din[7] 0.01fF
C1483 SA_OUT[7] PRE_A 0.00fF
C1484 PRE_CLSA ADC6_OUT[2] 0.09fF
C1485 Iref0 ADC4_OUT[1] 0.00fF
C1486 ADC6_OUT[0] Iref1 0.02fF
C1487 ADC1_OUT[1] ADC2_OUT[1] 0.01fF
C1488 VCLP ADC6_OUT[1] 0.91fF
C1489 ADC2_OUT[0] ADC3_OUT[2] 0.00fF
C1490 SAEN ADC5_OUT[1] 0.04fF
C1491 VDD ADC4_OUT[1] 1.58fF
C1492 a_5632_n6430# ADC9_OUT[0] 0.01fF
C1493 WWLD[0] WWLD[1] 0.86fF
C1494 ADC8_OUT[0] ADC8_OUT[2] 0.03fF
C1495 Din[1] PRE_A 0.00fF
C1496 Din[0] EN 0.01fF
C1497 PRE_SRAM WWLD[2] 0.00fF
C1498 VDD WWLD[3] 0.70fF
C1499 Din[8] Din[9] 0.02fF
C1500 a_5743_n6391# ADC7_OUT[1] 0.00fF
C1501 VCLP Iref3 0.14fF
C1502 WWLD[3] RWLB[1] 0.01fF
C1503 Din[12] PRE_A 0.00fF
C1504 VDD RWL[3] 2.83fF
C1505 WWL[0] RWL[1] 0.02fF
C1506 Din[11] EN 0.02fF
C1507 RWL[0] WWL[1] 0.01fF
C1508 m1_9142_5034# PRE_SRAM 0.14fF
C1509 ADC8_OUT[2] Iref2 0.02fF
C1510 ADC8_OUT[1] Iref3 0.01fF
C1511 ADC3_OUT[2] ADC4_OUT[3] 0.01fF
C1512 PRE_CLSA ADC2_OUT[0] 0.11fF
C1513 WWL[2] WWL[3] 0.10fF
C1514 RWL[1] RWLB[3] 0.01fF
C1515 PRE_A ADC4_OUT[0] 0.00fF
C1516 RWLB[1] RWL[3] 0.01fF
C1517 EN ADC3_OUT[0] 0.00fF
C1518 RWL[2] RWLB[2] 0.08fF
C1519 VDD WWL[7] 0.69fF
C1520 ADC0_OUT[0] ADC1_OUT[0] 0.01fF
C1521 WWL[1] WWL[4] 0.01fF
C1522 ADC14_OUT[2] ADC15_OUT[3] 0.02fF
C1523 ADC13_OUT[2] Iref3 0.01fF
C1524 Iref2 ADC13_OUT[3] 0.00fF
C1525 ADC9_OUT[2] ADC9_OUT[3] 1.32fF
C1526 RWLB[3] WWL[5] 0.02fF
C1527 VDD RWLB[10] 2.06fF
C1528 RWL[3] RWL[5] 0.02fF
C1529 WWL[3] RWLB[5] 0.01fF
C1530 WWL[4] RWLB[4] 21.69fF
C1531 a_5743_n6391# ADC14_OUT[0] 0.02fF
C1532 ADC11_OUT[3] ADC12_OUT[3] 0.02fF
C1533 a_5632_n6430# ADC11_OUT[1] 0.01fF
C1534 WWL[5] RWL[7] 0.01fF
C1535 RWLB[5] RWLB[6] 0.09fF
C1536 VDD RWL[14] 2.83fF
C1537 RWLB[4] RWLB[7] 0.00fF
C1538 RWL[5] WWL[7] 0.01fF
C1539 WWL[6] RWL[6] 22.38fF
C1540 SAEN ADC14_OUT[3] 0.02fF
C1541 ADC2_OUT[1] Iref1 0.01fF
C1542 PRE_CLSA ADC4_OUT[3] 0.10fF
C1543 ADC4_OUT[0] Iref2 0.01fF
C1544 SAEN ADC3_OUT[2] 0.04fF
C1545 ADC1_OUT[0] ADC2_OUT[3] 0.00fF
C1546 ADC0_OUT[1] ADC1_OUT[2] 0.01fF
C1547 VCLP ADC4_OUT[2] 0.95fF
C1548 m1_2819_5034# VDD 0.06fF
C1549 ADC12_OUT[0] VCLP 0.87fF
C1550 WWL[7] WWL[9] 0.03fF
C1551 RWLB[7] RWL[8] 1.23fF
C1552 RWL[6] RWLB[9] 0.00fF
C1553 VDD SA_OUT[1] 1.97fF
C1554 a_5743_n6391# ADC11_OUT[2] 0.92fF
C1555 RWLB[6] RWL[9] 0.01fF
C1556 RWL[7] RWLB[8] 0.01fF
C1557 VDD ADC2_OUT[2] 1.52fF
C1558 ADC6_OUT[1] ADC6_OUT[2] 3.84fF
C1559 ADC7_OUT[0] ADC7_OUT[3] 0.03fF
C1560 RWLB[9] WWL[10] 0.02fF
C1561 RWL[8] RWL[11] 0.00fF
C1562 PRE_CLSA ADC15_OUT[2] 0.07fF
C1563 VDD SA_OUT[12] 1.30fF
C1564 WWL[9] RWLB[10] 0.01fF
C1565 RWL[9] RWL[10] 0.09fF
C1566 WWL[8] RWLB[11] 0.00fF
C1567 VCLP ADC15_OUT[1] 0.76fF
C1568 ADC15_OUT[0] Iref1 0.02fF
C1569 RWLB[8] WWL[11] 0.01fF
C1570 WWL[0] Din[0] 0.00fF
C1571 PRE_SRAM Din[5] 0.01fF
C1572 WWLD[3] Din[1] 0.00fF
C1573 RWL[10] WWL[13] 0.00fF
C1574 WWL[11] RWL[12] 0.03fF
C1575 WWLD[2] Din[2] 0.00fF
C1576 RWL[11] WWL[12] 0.01fF
C1577 WWL[10] RWL[13] 0.00fF
C1578 WWLD[1] Din[3] 0.00fF
C1579 RWLB[10] RWLB[12] 0.02fF
C1580 WWLD[0] Din[4] 0.00fF
C1581 ADC12_OUT[0] ADC13_OUT[2] 0.00fF
C1582 VDD Din[6] 0.29fF
C1583 ADC6_OUT[2] Iref3 0.01fF
C1584 Iref2 ADC6_OUT[3] 0.00fF
C1585 ADC2_OUT[3] ADC3_OUT[3] 0.02fF
C1586 ADC0_OUT[0] VCLP 0.91fF
C1587 PRE_CLSA SAEN 0.27fF
C1588 ADC12_OUT[1] Iref2 0.01fF
C1589 ADC14_OUT[1] ADC14_OUT[2] 3.82fF
C1590 RWL[1] Din[7] 0.00fF
C1591 WWLD[1] Din[14] 0.00fF
C1592 WWL[1] Din[8] 0.00fF
C1593 RWLB[2] Din[3] 0.01fF
C1594 VDD EN 1.96fF
C1595 RWL[3] Din[1] 0.01fF
C1596 WWL[2] Din[5] 0.00fF
C1597 WWL[0] Din[11] 0.00fF
C1598 WWLD[2] Din[13] 0.00fF
C1599 WWLD[3] Din[12] 0.00fF
C1600 RWLB[0] Din[9] 0.01fF
C1601 RWL[12] RWLB[14] 0.01fF
C1602 RWL[13] RWLB[13] 0.08fF
C1603 WWL[12] WWL[15] 0.01fF
C1604 WWLD[0] Din[15] 0.00fF
C1605 RWLB[12] RWL[14] 0.01fF
C1606 RWL[2] Din[4] 0.00fF
C1607 RWLB[3] Din[0] 0.00fF
C1608 WWL[13] WWL[14] 0.10fF
C1609 RWLB[1] Din[6] 0.01fF
C1610 RWL[0] Din[10] 0.00fF
C1611 WWL[3] Din[2] 0.00fF
C1612 VDD ADC12_OUT[3] 1.58fF
C1613 m1_1670_5034# PRE_SRAM 0.14fF
C1614 ADC9_OUT[0] Iref0 0.03fF
C1615 PRE_CLSA ADC9_OUT[1] 0.10fF
C1616 m1_2819_5034# m1_3393_5034# 0.00fF
C1617 ADC10_OUT[0] SAEN 0.06fF
C1618 ADC4_OUT[0] ADC4_OUT[1] 5.48fF
C1619 ADC11_OUT[1] ADC11_OUT[3] 0.01fF
C1620 VDD ADC9_OUT[0] 2.27fF
C1621 RWL[14] WWLD[5] 0.00fF
C1622 RWLB[14] WWLD[4] 0.02fF
C1623 RWL[4] Din[9] 0.00fF
C1624 WWL[7] Din[1] 0.00fF
C1625 RWL[2] Din[15] 0.00fF
C1626 RWL[3] Din[12] 0.00fF
C1627 RWLB[6] Din[2] 0.01fF
C1628 RWLB[5] Din[5] 0.01fF
C1629 RWLB[2] Din[14] 0.01fF
C1630 RWL[5] Din[6] 0.00fF
C1631 RWL[7] Din[0] 0.00fF
C1632 WWL[15] RWLB[15] 21.69fF
C1633 RWL[6] Din[3] 0.00fF
C1634 RWLB[4] Din[8] 0.01fF
C1635 WWL[5] Din[7] 0.00fF
C1636 WWL[3] Din[13] 0.00fF
C1637 WWL[4] Din[10] 0.00fF
C1638 RWLB[3] Din[11] 0.01fF
C1639 WWL[6] Din[4] 0.00fF
C1640 SAEN ADC13_OUT[1] 0.03fF
C1641 ADC9_OUT[0] ADC10_OUT[1] 0.00fF
C1642 WWL[10] Din[3] 0.00fF
C1643 RWL[10] Din[2] 0.00fF
C1644 RWL[6] Din[14] 0.00fF
C1645 WWLD[7] PRE_VLSA 0.03fF
C1646 RWLB[9] Din[4] 0.01fF
C1647 RWL[9] Din[5] 0.00fF
C1648 RWL[8] Din[8] 0.00fF
C1649 WWLD[6] SA_OUT[0] 0.06fF
C1650 WWL[7] Din[12] 0.00fF
C1651 WWL[11] Din[0] 0.00fF
C1652 RWLB[7] Din[10] 0.01fF
C1653 RWLB[6] Din[13] 0.01fF
C1654 WWLD[5] SA_OUT[1] 0.04fF
C1655 RWLB[8] Din[7] 0.01fF
C1656 WWL[6] Din[15] 0.00fF
C1657 WWL[9] Din[6] 0.00fF
C1658 WWL[8] Din[9] 0.00fF
C1659 WWLD[4] SA_OUT[2] 0.01fF
C1660 RWLB[10] Din[1] 0.01fF
C1661 RWL[7] Din[11] 0.00fF
C1662 ADC0_OUT[1] Iref2 0.01fF
C1663 ADC2_OUT[0] Iref3 0.01fF
C1664 VCLP ADC2_OUT[3] 1.02fF
C1665 SAEN ADC1_OUT[3] 0.02fF
C1666 VDD ADC0_OUT[3] 1.55fF
C1667 m1_3393_5034# Din[6] 0.00fF
C1668 RWLB[9] Din[15] 0.01fF
C1669 WWLD[5] SA_OUT[12] 0.00fF
C1670 SA_OUT[1] SA_OUT[7] 0.00fF
C1671 RWL[10] Din[13] 0.00fF
C1672 RWL[11] Din[10] 0.00fF
C1673 WWL[13] Din[5] 0.00fF
C1674 RWLB[10] Din[12] 0.01fF
C1675 RWL[12] Din[7] 0.01fF
C1676 SA_OUT[0] SA_OUT[8] 0.00fF
C1677 SA_OUT[3] SA_OUT[5] 0.01fF
C1678 WWLD[6] SA_OUT[11] 0.00fF
C1679 RWLB[12] Din[6] 0.01fF
C1680 WWLD[7] SA_OUT[10] 0.02fF
C1681 SA_OUT[2] SA_OUT[6] 0.01fF
C1682 WWL[10] Din[14] 0.00fF
C1683 WWL[14] Din[2] 0.00fF
C1684 WWL[12] Din[8] 0.00fF
C1685 RWL[13] Din[4] 0.00fF
C1686 RWLB[14] Din[0] 0.00fF
C1687 PRE_VLSA SA_OUT[9] 0.27fF
C1688 RWL[14] Din[1] 0.00fF
C1689 WWL[11] Din[11] 0.00fF
C1690 RWLB[11] Din[9] 0.01fF
C1691 RWLB[13] Din[3] 0.01fF
C1692 ADC5_OUT[1] ADC5_OUT[3] 0.01fF
C1693 SA_OUT[9] SA_OUT[10] 4.06fF
C1694 WWLD[6] Din[5] 0.00fF
C1695 SA_OUT[8] SA_OUT[11] 0.02fF
C1696 RWLB[14] Din[11] 0.01fF
C1697 RWL[14] Din[12] 0.00fF
C1698 SA_OUT[6] SA_OUT[13] 0.03fF
C1699 WWL[15] Din[10] 0.00fF
C1700 SA_OUT[0] Din[2] 0.02fF
C1701 RWLB[13] Din[14] 0.01fF
C1702 SA_OUT[1] Din[1] 0.00fF
C1703 SA_OUT[3] WE 0.01fF
C1704 RWL[13] Din[15] 0.00fF
C1705 WWL[14] Din[13] 0.00fF
C1706 SA_OUT[7] SA_OUT[12] 0.02fF
C1707 PRE_VLSA Din[3] 0.02fF
C1708 RWLB[15] Din[8] 0.01fF
C1709 WWLD[7] Din[4] 0.00fF
C1710 SA_OUT[4] SA_OUT[15] 0.01fF
C1711 WWLD[5] Din[6] 0.00fF
C1712 SA_OUT[5] SA_OUT[14] 0.01fF
C1713 RWL[15] Din[9] 0.00fF
C1714 WWLD[4] Din[7] 0.00fF
C1715 m1_7993_5034# Din[14] 0.00fF
C1716 ADC4_OUT[3] Iref3 0.01fF
C1717 Iref0 ADC11_OUT[1] 0.00fF
C1718 PRE_VLSA Din[14] 0.02fF
C1719 SA_OUT[4] Din[9] 0.01fF
C1720 SA_OUT[5] Din[8] 0.01fF
C1721 SA_OUT[3] Din[10] 0.01fF
C1722 SA_OUT[0] Din[13] 0.02fF
C1723 SA_OUT[6] Din[7] 0.01fF
C1724 WWLD[7] Din[15] 0.00fF
C1725 SA_OUT[1] Din[12] 0.01fF
C1726 SA_OUT[2] Din[11] 0.01fF
C1727 SA_OUT[14] WE 0.02fF
C1728 VDD ADC11_OUT[1] 1.57fF
C1729 a_5632_n6430# PRE_CLSA 0.03fF
C1730 ADC10_OUT[1] ADC11_OUT[1] 0.01fF
C1731 SA_OUT[12] Din[12] 0.00fF
C1732 SA_OUT[9] Din[15] 0.01fF
C1733 Din[3] Din[4] 0.02fF
C1734 SA_OUT[11] Din[13] 0.01fF
C1735 SA_OUT[10] Din[14] 0.01fF
C1736 WE Din[8] 0.01fF
C1737 SA_OUT[7] EN 0.00fF
C1738 SA_OUT[8] PRE_A 0.00fF
C1739 Iref0 ADC5_OUT[1] 0.00fF
C1740 SAEN ADC6_OUT[1] 0.04fF
C1741 Iref2 ADC15_OUT[3] 0.01fF
C1742 ADC7_OUT[0] Iref1 0.02fF
C1743 PRE_CLSA ADC7_OUT[2] 0.09fF
C1744 ADC15_OUT[2] Iref3 0.01fF
C1745 ADC3_OUT[0] ADC3_OUT[2] 0.03fF
C1746 VCLP ADC7_OUT[1] 0.90fF
C1747 a_5632_n6430# ADC10_OUT[0] 0.01fF
C1748 a_5743_n6391# VCLP 0.12fF
C1749 VDD ADC5_OUT[1] 1.57fF
C1750 WWLD[0] WWLD[2] 0.03fF
C1751 VDD WWL[0] 0.69fF
C1752 Din[1] EN 0.02fF
C1753 Din[2] PRE_A 0.00fF
C1754 ADC8_OUT[0] ADC9_OUT[2] 0.00fF
C1755 ADC7_OUT[1] ADC8_OUT[1] 0.01fF
C1756 ADC12_OUT[3] ADC13_OUT[3] 0.02fF
C1757 m1_1670_5034# Din[2] 0.00fF
C1758 a_5632_n6430# ADC13_OUT[1] 0.01fF
C1759 PRE_A ADC11_OUT[0] 0.00fF
C1760 SAEN Iref3 0.16fF
C1761 a_5743_n6391# ADC8_OUT[1] 0.01fF
C1762 Din[13] PRE_A 0.00fF
C1763 Din[12] EN 0.00fF
C1764 RWL[0] RWL[1] 0.09fF
C1765 WWLD[3] WWL[2] 0.01fF
C1766 Din[14] Din[15] 0.02fF
C1767 VDD RWLB[3] 2.06fF
C1768 WWL[0] RWLB[1] 0.01fF
C1769 RWLB[0] WWL[1] 0.02fF
C1770 m1_3968_5034# VDD 0.06fF
C1771 ADC14_OUT[0] VCLP 0.87fF
C1772 a_5743_n6391# ADC13_OUT[2] 0.96fF
C1773 ADC9_OUT[2] Iref2 0.02fF
C1774 ADC4_OUT[2] ADC4_OUT[3] 1.29fF
C1775 ADC9_OUT[1] Iref3 0.01fF
C1776 RWL[2] WWL[3] 0.01fF
C1777 EN ADC4_OUT[0] 0.00fF
C1778 PRE_CLSA ADC3_OUT[0] 0.11fF
C1779 WWL[2] RWL[3] 0.02fF
C1780 RWL[1] WWL[4] 0.00fF
C1781 RWLB[1] RWLB[3] 0.02fF
C1782 VDD RWL[7] 2.83fF
C1783 PRE_A ADC5_OUT[0] 0.00fF
C1784 WWL[1] RWL[4] 0.01fF
C1785 m1_6269_5033# Din[10] 0.00fF
C1786 ADC9_OUT[2] ADC10_OUT[3] 0.01fF
C1787 WWL[4] WWL[5] 0.10fF
C1788 ADC6_OUT[0] ADC7_OUT[0] 0.01fF
C1789 RWL[4] RWLB[4] 0.08fF
C1790 RWLB[3] RWL[5] 0.01fF
C1791 WWL[3] WWL[6] 0.01fF
C1792 VDD WWL[11] 0.70fF
C1793 RWL[3] RWLB[5] 0.01fF
C1794 ADC13_OUT[0] ADC14_OUT[2] 0.00fF
C1795 PRE_CLSA ADC11_OUT[3] 0.10fF
C1796 ADC11_OUT[0] Iref2 0.01fF
C1797 VCLP ADC11_OUT[2] 0.02fF
C1798 WWL[6] RWLB[6] 21.69fF
C1799 RWL[5] RWL[7] 0.02fF
C1800 RWLB[5] WWL[7] 0.02fF
C1801 VDD RWLB[14] 2.06fF
C1802 WWL[5] RWLB[7] 0.01fF
C1803 ADC15_OUT[1] ADC15_OUT[2] 3.83fF
C1804 ADC14_OUT[1] Iref2 0.01fF
C1805 ADC10_OUT[0] ADC11_OUT[3] 0.00fF
C1806 ADC3_OUT[1] Iref1 0.01fF
C1807 ADC5_OUT[0] Iref2 0.01fF
C1808 ADC2_OUT[0] ADC2_OUT[3] 0.03fF
C1809 SAEN ADC4_OUT[2] 0.04fF
C1810 PRE_CLSA ADC5_OUT[3] 0.10fF
C1811 ADC1_OUT[1] ADC1_OUT[2] 3.82fF
C1812 VDD ADC14_OUT[3] 1.63fF
C1813 VCLP ADC5_OUT[2] 0.94fF
C1814 WWL[7] RWL[9] 0.01fF
C1815 VDD SA_OUT[2] 1.84fF
C1816 RWLB[6] RWLB[9] 0.00fF
C1817 WWL[8] RWL[8] 22.38fF
C1818 RWL[7] WWL[9] 0.01fF
C1819 RWLB[7] RWLB[8] 0.09fF
C1820 m1_2819_5034# PRE_SRAM 0.14fF
C1821 VDD ADC3_OUT[2] 1.53fF
C1822 m1_3393_5034# m1_3968_5034# 0.00fF
C1823 ADC12_OUT[0] SAEN 0.06fF
C1824 ADC12_OUT[1] ADC12_OUT[3] 0.01fF
C1825 ADC6_OUT[1] ADC7_OUT[2] 0.01fF
C1826 ADC7_OUT[0] ADC8_OUT[3] 0.00fF
C1827 SAEN ADC15_OUT[1] 0.02fF
C1828 VDD SA_OUT[13] 1.33fF
C1829 RWLB[8] RWL[11] 0.01fF
C1830 WWL[9] WWL[11] 0.03fF
C1831 RWL[8] RWLB[11] 0.00fF
C1832 RWLB[9] RWL[10] 1.23fF
C1833 RWL[9] RWLB[10] 0.01fF
C1834 WWLD[2] Din[3] 0.00fF
C1835 WWLD[0] Din[5] 0.00fF
C1836 PRE_SRAM Din[6] 0.01fF
C1837 VDD Din[7] 0.26fF
C1838 RWL[10] RWL[13] 0.00fF
C1839 WWL[0] Din[1] 0.00fF
C1840 RWL[0] Din[0] 0.00fF
C1841 WWLD[1] Din[4] 0.00fF
C1842 RWL[11] RWL[12] 0.08fF
C1843 RWLB[10] WWL[13] 0.00fF
C1844 a_5632_n6430# Iref3 0.00fF
C1845 RWLB[11] WWL[12] 0.02fF
C1846 WWL[11] RWLB[12] 0.01fF
C1847 WWLD[3] Din[2] 0.00fF
C1848 WWL[10] RWLB[13] 0.00fF
C1849 Iref2 ADC7_OUT[3] 0.00fF
C1850 ADC7_OUT[2] Iref3 0.01fF
C1851 ADC0_OUT[0] SAEN 0.08fF
C1852 PRE_CLSA Iref0 0.01fF
C1853 ADC1_OUT[0] VCLP 0.90fF
C1854 RWLB[12] RWLB[14] 0.02fF
C1855 RWL[2] Din[5] 0.00fF
C1856 RWLB[1] Din[7] 0.01fF
C1857 RWLB[3] Din[1] 0.01fF
C1858 RWLB[2] Din[4] 0.01fF
C1859 WWLD[1] Din[15] 0.00fF
C1860 WWL[2] Din[6] 0.00fF
C1861 WWLD[2] Din[14] 0.00fF
C1862 RWL[1] Din[8] 0.00fF
C1863 WWL[12] RWL[15] 0.01fF
C1864 WWL[3] Din[3] 0.00fF
C1865 WWL[13] RWL[14] 0.02fF
C1866 RWL[13] WWL[14] 0.01fF
C1867 RWL[12] WWL[15] 0.00fF
C1868 WWL[4] Din[0] 0.00fF
C1869 VDD PRE_CLSA 31.52fF
C1870 WWL[1] Din[9] 0.00fF
C1871 WWL[0] Din[12] 0.00fF
C1872 RWL[3] Din[2] 0.00fF
C1873 RWLB[0] Din[10] 0.01fF
C1874 WWLD[3] Din[13] 0.00fF
C1875 RWL[0] Din[11] 0.00fF
C1876 ADC8_OUT[3] ADC9_OUT[3] 0.02fF
C1877 ADC4_OUT[0] ADC5_OUT[1] 0.00fF
C1878 ADC10_OUT[0] Iref0 0.03fF
C1879 PRE_CLSA ADC10_OUT[1] 0.10fF
C1880 RWL[3] Din[13] 0.00fF
C1881 WWL[3] Din[14] 0.00fF
C1882 RWLB[2] Din[15] 0.01fF
C1883 WWL[4] Din[11] 0.00fF
C1884 RWL[5] Din[7] 0.00fF
C1885 RWL[7] Din[1] 0.00fF
C1886 RWLB[6] Din[3] 0.01fF
C1887 RWLB[7] Din[0] 0.00fF
C1888 VDD ADC10_OUT[0] 2.28fF
C1889 WWL[15] WWLD[4] 0.10fF
C1890 WWL[5] Din[8] 0.00fF
C1891 RWLB[3] Din[12] 0.01fF
C1892 RWLB[14] WWLD[5] 0.01fF
C1893 RWLB[4] Din[9] 0.01fF
C1894 WWL[6] Din[5] 0.00fF
C1895 RWL[4] Din[10] 0.00fF
C1896 RWL[15] RWLB[15] 0.08fF
C1897 RWL[6] Din[4] 0.00fF
C1898 RWLB[5] Din[6] 0.01fF
C1899 WWL[7] Din[2] 0.00fF
C1900 Iref0 ADC13_OUT[1] 0.00fF
C1901 ADC10_OUT[0] ADC10_OUT[1] 5.53fF
C1902 VDD ADC13_OUT[1] 1.58fF
C1903 WWL[7] Din[13] 0.00fF
C1904 WWL[10] Din[4] 0.00fF
C1905 WWLD[6] SA_OUT[1] 0.18fF
C1906 WWL[11] Din[1] 0.00fF
C1907 WWLD[5] SA_OUT[2] 0.03fF
C1908 WWL[9] Din[7] 0.00fF
C1909 RWLB[8] Din[8] 0.01fF
C1910 WWL[8] Din[10] 0.00fF
C1911 RWL[9] Din[6] 0.00fF
C1912 WWLD[4] SA_OUT[3] 0.00fF
C1913 RWL[7] Din[12] 0.00fF
C1914 WWLD[7] SA_OUT[0] 0.06fF
C1915 RWL[6] Din[15] 0.00fF
C1916 RWLB[10] Din[2] 0.01fF
C1917 RWLB[7] Din[11] 0.01fF
C1918 RWLB[6] Din[14] 0.01fF
C1919 RWLB[9] Din[5] 0.01fF
C1920 RWL[10] Din[3] 0.00fF
C1921 RWL[11] Din[0] 0.00fF
C1922 RWL[8] Din[9] 0.00fF
C1923 SAEN ADC2_OUT[3] 0.02fF
C1924 VCLP ADC3_OUT[3] 1.03fF
C1925 ADC1_OUT[1] Iref2 0.01fF
C1926 ADC0_OUT[1] ADC0_OUT[3] 0.01fF
C1927 ADC3_OUT[0] Iref3 0.01fF
C1928 ADC11_OUT[1] ADC12_OUT[1] 0.01fF
C1929 VDD ADC1_OUT[3] 1.58fF
C1930 SA_OUT[3] SA_OUT[6] 0.01fF
C1931 RWLB[13] Din[4] 0.01fF
C1932 SA_OUT[0] SA_OUT[9] 0.00fF
C1933 RWL[13] Din[5] 0.00fF
C1934 WWL[14] Din[3] 0.00fF
C1935 WWL[12] Din[9] 0.00fF
C1936 RWL[10] Din[14] 0.00fF
C1937 RWL[11] Din[11] 0.00fF
C1938 RWLB[14] Din[1] 0.01fF
C1939 WWL[13] Din[6] 0.00fF
C1940 WWL[11] Din[12] 0.00fF
C1941 WWLD[7] SA_OUT[11] 0.02fF
C1942 PRE_VLSA SA_OUT[10] 0.25fF
C1943 RWLB[11] Din[10] 0.01fF
C1944 RWL[14] Din[2] 0.00fF
C1945 SA_OUT[4] SA_OUT[5] 3.39fF
C1946 WWLD[6] SA_OUT[12] 0.00fF
C1947 RWLB[10] Din[13] 0.01fF
C1948 SA_OUT[2] SA_OUT[7] 0.01fF
C1949 RWLB[12] Din[7] 0.01fF
C1950 RWL[12] Din[8] 0.00fF
C1951 WWLD[5] SA_OUT[13] 0.00fF
C1952 WWL[10] Din[15] 0.00fF
C1953 SA_OUT[1] SA_OUT[8] 0.00fF
C1954 WWL[15] Din[0] 0.00fF
C1955 a_5632_n6430# ADC12_OUT[0] 0.01fF
C1956 ADC5_OUT[2] ADC6_OUT[2] 0.01fF
C1957 ADC5_OUT[1] ADC6_OUT[3] 0.00fF
C1958 ADC13_OUT[3] ADC14_OUT[3] 0.02fF
C1959 ADC11_OUT[3] Iref3 0.01fF
C1960 SA_OUT[9] SA_OUT[11] 0.02fF
C1961 SA_OUT[0] Din[3] 0.02fF
C1962 SA_OUT[1] Din[2] 0.01fF
C1963 WWLD[5] Din[7] 0.00fF
C1964 WWLD[7] Din[5] 0.00fF
C1965 WWLD[6] Din[6] 0.00fF
C1966 RWL[15] Din[10] 0.00fF
C1967 WWL[15] Din[11] 0.00fF
C1968 RWLB[15] Din[9] 0.01fF
C1969 WWLD[4] Din[8] 0.00fF
C1970 SA_OUT[7] SA_OUT[13] 0.02fF
C1971 SA_OUT[8] SA_OUT[12] 0.02fF
C1972 SA_OUT[5] SA_OUT[15] 0.02fF
C1973 SA_OUT[6] SA_OUT[14] 0.04fF
C1974 RWLB[14] Din[12] 0.01fF
C1975 RWL[14] Din[13] 0.00fF
C1976 WWL[14] Din[14] 0.00fF
C1977 PRE_VLSA Din[4] 0.02fF
C1978 SA_OUT[4] WE 0.01fF
C1979 RWLB[13] Din[15] 0.01fF
C1980 a_5632_n6430# ADC15_OUT[1] 0.00fF
C1981 SA_OUT[6] Din[8] 0.01fF
C1982 ADC5_OUT[3] Iref3 0.01fF
C1983 SA_OUT[1] Din[13] 0.01fF
C1984 SA_OUT[2] Din[12] 0.01fF
C1985 m1_5118_5034# VDD 0.06fF
C1986 SA_OUT[3] Din[11] 0.01fF
C1987 SA_OUT[0] Din[14] 0.02fF
C1988 PRE_VLSA Din[15] 0.02fF
C1989 SA_OUT[4] Din[10] 0.01fF
C1990 SA_OUT[7] Din[7] 0.00fF
C1991 SA_OUT[15] WE 0.01fF
C1992 SA_OUT[5] Din[9] 0.01fF
C1993 a_5743_n6391# ADC15_OUT[2] 0.74fF
C1994 WE Din[9] 0.01fF
C1995 VCLP ADC8_OUT[1] 0.92fF
C1996 SA_OUT[11] Din[14] 0.01fF
C1997 SAEN ADC7_OUT[1] 0.03fF
C1998 Iref0 ADC6_OUT[1] 0.00fF
C1999 ADC3_OUT[0] ADC4_OUT[2] 0.00fF
C2000 SA_OUT[8] EN 0.00fF
C2001 ADC2_OUT[1] ADC3_OUT[1] 0.01fF
C2002 SA_OUT[12] Din[13] 0.01fF
C2003 ADC8_OUT[0] Iref1 0.02fF
C2004 PRE_CLSA ADC8_OUT[2] 0.09fF
C2005 SA_OUT[10] Din[15] 0.01fF
C2006 SA_OUT[9] PRE_A 0.00fF
C2007 VDD ADC6_OUT[1] 1.56fF
C2008 a_5743_n6391# SAEN 0.00fF
C2009 ADC13_OUT[0] Iref2 0.01fF
C2010 PRE_CLSA ADC13_OUT[3] 0.10fF
C2011 WWLD[0] WWLD[3] 0.01fF
C2012 VDD RWL[0] 2.83fF
C2013 Din[2] EN 0.00fF
C2014 WWLD[1] WWLD[2] 0.70fF
C2015 Din[3] PRE_A 0.00fF
C2016 ADC15_OUT[0] ADC14_OUT[2] 0.00fF
C2017 ADC14_OUT[0] ADC15_OUT[2] 0.00fF
C2018 Din[9] Din[10] 0.02fF
C2019 VCLP ADC13_OUT[2] 0.02fF
C2020 ADC9_OUT[0] ADC9_OUT[2] 0.03fF
C2021 m1_1670_5034# Din[3] 0.00fF
C2022 a_5743_n6391# ADC9_OUT[1] 0.01fF
C2023 Iref0 Iref3 0.01fF
C2024 Iref1 Iref2 1.96fF
C2025 WWLD[3] RWL[2] 0.01fF
C2026 Din[14] PRE_A 0.00fF
C2027 RWLB[0] RWL[1] 1.23fF
C2028 RWL[0] RWLB[1] 0.01fF
C2029 WWL[0] WWL[2] 0.03fF
C2030 Din[13] EN 0.02fF
C2031 VDD WWL[4] 0.70fF
C2032 ADC11_OUT[0] ADC12_OUT[3] 0.00fF
C2033 VDD Iref3 0.41fF
C2034 m1_3968_5034# PRE_SRAM 0.14fF
C2035 m1_3968_5034# m1_4543_5034# 0.00fF
C2036 ADC14_OUT[0] SAEN 0.06fF
C2037 ADC4_OUT[2] ADC5_OUT[3] 0.01fF
C2038 ADC10_OUT[1] Iref3 0.01fF
C2039 ADC13_OUT[1] ADC13_OUT[3] 0.01fF
C2040 ADC10_OUT[2] Iref2 0.02fF
C2041 RWL[2] RWL[3] 0.09fF
C2042 RWL[1] RWL[4] 0.00fF
C2043 EN ADC5_OUT[0] 0.00fF
C2044 VDD RWLB[7] 2.06fF
C2045 WWL[2] RWLB[3] 0.01fF
C2046 RWLB[1] WWL[4] 0.00fF
C2047 PRE_CLSA ADC4_OUT[0] 0.11fF
C2048 RWLB[2] WWL[3] 0.02fF
C2049 ADC1_OUT[0] ADC2_OUT[0] 0.01fF
C2050 WWL[1] RWLB[4] 0.00fF
C2051 PRE_A ADC6_OUT[0] 0.00fF
C2052 m1_6269_5033# Din[11] 0.00fF
C2053 ADC10_OUT[2] ADC10_OUT[3] 1.34fF
C2054 RWL[4] WWL[5] 0.01fF
C2055 WWL[3] RWL[6] 0.00fF
C2056 RWL[3] WWL[6] 0.00fF
C2057 WWL[4] RWL[5] 0.02fF
C2058 RWLB[3] RWLB[5] 0.02fF
C2059 VDD RWL[11] 2.83fF
C2060 SAEN ADC11_OUT[2] 0.01fF
C2061 RWL[5] RWLB[7] 0.01fF
C2062 RWLB[5] RWL[7] 0.01fF
C2063 WWL[6] WWL[7] 0.10fF
C2064 WWL[5] WWL[8] 0.01fF
C2065 RWL[6] RWLB[6] 0.08fF
C2066 VDD WWL[15] 0.69fF
C2067 VCLP ADC6_OUT[2] 0.93fF
C2068 PRE_CLSA ADC6_OUT[3] 0.10fF
C2069 ADC4_OUT[1] Iref1 0.01fF
C2070 SAEN ADC5_OUT[2] 0.04fF
C2071 ADC1_OUT[1] ADC2_OUT[2] 0.01fF
C2072 ADC6_OUT[0] Iref2 0.01fF
C2073 ADC2_OUT[0] ADC3_OUT[3] 0.00fF
C2074 RWL[7] RWL[9] 0.02fF
C2075 RWLB[7] WWL[9] 0.02fF
C2076 WWL[8] RWLB[8] 21.69fF
C2077 WWL[7] RWLB[9] 0.01fF
C2078 VDD SA_OUT[3] 1.73fF
C2079 PRE_CLSA ADC12_OUT[1] 0.10fF
C2080 VDD ADC4_OUT[2] 1.52fF
C2081 ADC12_OUT[0] Iref0 0.03fF
C2082 a_5632_n6430# ADC7_OUT[1] 0.01fF
C2083 VDD ADC12_OUT[0] 2.27fF
C2084 ADC8_OUT[0] ADC8_OUT[3] 0.03fF
C2085 ADC7_OUT[1] ADC7_OUT[2] 3.85fF
C2086 a_5743_n6391# a_5632_n6430# 14.25fF
C2087 RWL[9] WWL[11] 0.01fF
C2088 Iref0 ADC15_OUT[1] 0.32fF
C2089 RWLB[9] RWLB[10] 0.09fF
C2090 VDD SA_OUT[14] 1.38fF
C2091 RWLB[8] RWLB[11] 0.00fF
C2092 WWL[10] RWL[10] 22.38fF
C2093 WWL[9] RWL[11] 0.01fF
C2094 ADC11_OUT[0] ADC11_OUT[1] 5.54fF
C2095 a_5743_n6391# ADC7_OUT[2] 0.16fF
C2096 VDD ADC15_OUT[1] 1.54fF
C2097 ADC12_OUT[1] ADC13_OUT[1] 0.01fF
C2098 WWL[11] WWL[13] 0.03fF
C2099 RWLB[11] RWL[12] 0.97fF
C2100 WWLD[1] Din[5] 0.00fF
C2101 WWLD[2] Din[4] 0.00fF
C2102 RWL[0] Din[1] 0.00fF
C2103 RWL[11] RWLB[12] 0.01fF
C2104 WWL[0] Din[2] 0.00fF
C2105 WWLD[0] Din[6] 0.00fF
C2106 WWLD[3] Din[3] 0.00fF
C2107 RWLB[0] Din[0] 0.00fF
C2108 PRE_SRAM Din[7] 0.01fF
C2109 RWLB[10] RWL[13] 0.01fF
C2110 VDD Din[8] 0.29fF
C2111 m1_4543_5034# Din[7] 0.00fF
C2112 ADC8_OUT[2] Iref3 0.01fF
C2113 Iref2 ADC8_OUT[3] 0.00fF
C2114 ADC3_OUT[3] ADC4_OUT[3] 0.02fF
C2115 ADC0_OUT[0] Iref0 0.02fF
C2116 ADC1_OUT[0] SAEN 0.07fF
C2117 PRE_CLSA ADC0_OUT[1] 0.11fF
C2118 ADC2_OUT[0] VCLP 0.88fF
C2119 a_5632_n6430# ADC14_OUT[0] 0.01fF
C2120 WWL[2] Din[7] 0.00fF
C2121 WWLD[2] Din[15] 0.00fF
C2122 WWLD[3] Din[14] 0.00fF
C2123 RWLB[0] Din[11] 0.01fF
C2124 RWLB[13] WWL[14] 0.02fF
C2125 WWL[13] RWLB[14] 0.01fF
C2126 WWL[12] RWLB[15] 0.00fF
C2127 WWL[1] Din[10] 0.00fF
C2128 RWLB[12] WWL[15] 0.01fF
C2129 RWL[1] Din[9] 0.00fF
C2130 RWL[2] Din[6] 0.00fF
C2131 WWL[0] Din[13] 0.00fF
C2132 WWL[4] Din[1] 0.00fF
C2133 RWL[0] Din[12] 0.00fF
C2134 RWL[4] Din[0] 0.00fF
C2135 RWL[3] Din[3] 0.00fF
C2136 WWL[3] Din[4] 0.00fF
C2137 RWLB[1] Din[8] 0.01fF
C2138 RWL[13] RWL[14] 0.09fF
C2139 RWLB[2] Din[5] 0.01fF
C2140 RWL[12] RWL[15] 0.00fF
C2141 RWLB[3] Din[2] 0.01fF
C2142 VDD ADC0_OUT[0] 2.27fF
C2143 ADC13_OUT[3] Iref3 0.01fF
C2144 ADC14_OUT[3] ADC15_OUT[3] 0.03fF
C2145 ADC5_OUT[0] ADC5_OUT[1] 5.50fF
C2146 RWLB[3] Din[13] 0.01fF
C2147 RWLB[4] Din[10] 0.01fF
C2148 WWL[8] Din[0] 0.00fF
C2149 RWL[3] Din[14] 0.00fF
C2150 WWL[5] Din[9] 0.00fF
C2151 RWLB[5] Din[7] 0.01fF
C2152 RWL[6] Din[5] 0.00fF
C2153 RWLB[6] Din[4] 0.01fF
C2154 RWL[15] WWLD[4] 0.01fF
C2155 WWL[3] Din[15] 0.00fF
C2156 WWL[4] Din[12] 0.00fF
C2157 RWL[5] Din[8] 0.00fF
C2158 WWL[7] Din[3] 0.00fF
C2159 WWL[6] Din[6] 0.00fF
C2160 WWL[15] WWLD[5] 0.03fF
C2161 RWL[4] Din[11] 0.00fF
C2162 RWL[7] Din[2] 0.00fF
C2163 RWLB[7] Din[1] 0.01fF
C2164 m1_9142_5034# Din[15] 0.00fF
C2165 m1_6269_5033# VDD 0.04fF
C2166 a_5632_n6430# ADC11_OUT[2] 0.02fF
C2167 RWLB[8] Din[9] 0.01fF
C2168 WWL[7] Din[14] 0.00fF
C2169 RWLB[7] Din[12] 0.01fF
C2170 RWLB[6] Din[15] 0.01fF
C2171 RWLB[11] Din[0] 0.00fF
C2172 WWLD[7] SA_OUT[1] 0.07fF
C2173 RWLB[10] Din[3] 0.01fF
C2174 RWL[8] Din[10] 0.00fF
C2175 WWL[8] Din[11] 0.00fF
C2176 RWL[11] Din[1] 0.01fF
C2177 PRE_VLSA SA_OUT[0] 0.12fF
C2178 WWL[10] Din[5] 0.00fF
C2179 WWLD[6] SA_OUT[2] 0.05fF
C2180 WWLD[5] SA_OUT[3] 0.02fF
C2181 WWL[11] Din[2] 0.00fF
C2182 RWL[10] Din[4] 0.00fF
C2183 WWL[9] Din[8] 0.00fF
C2184 RWL[9] Din[7] 0.00fF
C2185 RWLB[9] Din[6] 0.01fF
C2186 RWL[7] Din[13] 0.00fF
C2187 ADC2_OUT[1] Iref2 0.01fF
C2188 ADC0_OUT[2] ADC1_OUT[2] 0.01fF
C2189 SAEN ADC3_OUT[3] 0.02fF
C2190 ADC0_OUT[1] ADC1_OUT[3] 0.00fF
C2191 VCLP ADC4_OUT[3] 1.03fF
C2192 ADC4_OUT[0] Iref3 0.01fF
C2193 VDD ADC2_OUT[3] 1.58fF
C2194 SA_OUT[1] SA_OUT[9] 0.00fF
C2195 RWLB[14] Din[2] 0.01fF
C2196 RWL[15] Din[0] 0.00fF
C2197 RWL[14] Din[3] 0.00fF
C2198 SA_OUT[3] SA_OUT[7] 0.01fF
C2199 RWLB[12] Din[8] 0.01fF
C2200 WWL[14] Din[4] 0.00fF
C2201 WWLD[5] SA_OUT[14] 0.00fF
C2202 SA_OUT[4] SA_OUT[6] 0.01fF
C2203 RWL[13] Din[6] 0.00fF
C2204 PRE_VLSA SA_OUT[11] 0.22fF
C2205 RWL[12] Din[9] 0.00fF
C2206 WWLD[6] SA_OUT[13] 0.00fF
C2207 SA_OUT[2] SA_OUT[8] 0.01fF
C2208 WWL[15] Din[1] 0.00fF
C2209 RWLB[11] Din[11] 0.01fF
C2210 RWLB[13] Din[5] 0.01fF
C2211 RWL[10] Din[15] 0.00fF
C2212 WWL[12] Din[10] 0.00fF
C2213 RWL[11] Din[12] 0.00fF
C2214 RWLB[10] Din[14] 0.01fF
C2215 WWLD[7] SA_OUT[12] 0.02fF
C2216 SA_OUT[0] SA_OUT[10] 0.00fF
C2217 WWL[13] Din[7] 0.00fF
C2218 WWL[11] Din[13] 0.00fF
C2219 ADC6_OUT[1] ADC6_OUT[3] 0.01fF
C2220 VCLP ADC15_OUT[2] 0.00fF
C2221 PRE_CLSA ADC15_OUT[3] 0.07fF
C2222 ADC15_OUT[0] Iref2 0.01fF
C2223 RWLB[14] Din[13] 0.01fF
C2224 WWLD[4] Din[9] 0.00fF
C2225 SA_OUT[0] Din[4] 0.02fF
C2226 WWL[14] Din[15] 0.00fF
C2227 PRE_VLSA Din[5] 0.02fF
C2228 SA_OUT[6] SA_OUT[15] 0.04fF
C2229 SA_OUT[8] SA_OUT[13] 0.02fF
C2230 RWL[15] Din[11] 0.00fF
C2231 WWLD[7] Din[6] 0.00fF
C2232 SA_OUT[9] SA_OUT[12] 0.02fF
C2233 SA_OUT[5] WE 0.01fF
C2234 SA_OUT[2] Din[2] 0.00fF
C2235 SA_OUT[10] SA_OUT[11] 3.89fF
C2236 RWL[14] Din[14] 0.00fF
C2237 WWLD[6] Din[7] 0.00fF
C2238 WWLD[5] Din[8] 0.00fF
C2239 SA_OUT[7] SA_OUT[14] 0.02fF
C2240 WWL[15] Din[12] 0.00fF
C2241 RWLB[15] Din[10] 0.01fF
C2242 SA_OUT[1] Din[3] 0.01fF
C2243 ADC12_OUT[0] ADC13_OUT[3] 0.00fF
C2244 SA_OUT[7] Din[8] 0.01fF
C2245 PRE_VLSA PRE_A 0.05fF
C2246 SA_OUT[1] Din[14] 0.01fF
C2247 SA_OUT[5] Din[10] 0.01fF
C2248 ADC6_OUT[3] Iref3 0.01fF
C2249 SA_OUT[6] Din[9] 0.01fF
C2250 m1_5118_5034# PRE_SRAM 0.14fF
C2251 SA_OUT[4] Din[11] 0.01fF
C2252 SA_OUT[2] Din[13] 0.01fF
C2253 SA_OUT[3] Din[12] 0.01fF
C2254 SA_OUT[0] Din[15] 0.02fF
C2255 m1_4543_5034# m1_5118_5034# 0.00fF
C2256 VCLP SAEN 103.73fF
C2257 ADC12_OUT[1] Iref3 0.01fF
C2258 ADC14_OUT[1] ADC14_OUT[3] 0.01fF
C2259 ADC12_OUT[2] Iref2 0.02fF
C2260 SA_OUT[13] Din[13] 0.00fF
C2261 SA_OUT[10] PRE_A 0.00fF
C2262 SA_OUT[9] EN 0.00fF
C2263 WE Din[10] 0.01fF
C2264 SA_OUT[12] Din[14] 0.01fF
C2265 Din[4] Din[5] 0.02fF
C2266 SA_OUT[11] Din[15] 0.01fF
C2267 ADC4_OUT[0] ADC4_OUT[2] 0.03fF
C2268 VCLP ADC9_OUT[1] 0.92fF
C2269 ADC9_OUT[0] Iref1 0.02fF
C2270 SAEN ADC8_OUT[1] 0.03fF
C2271 Iref0 ADC7_OUT[1] 0.00fF
C2272 PRE_CLSA ADC9_OUT[2] 0.09fF
C2273 ADC11_OUT[2] ADC11_OUT[3] 1.35fF
C2274 VDD ADC7_OUT[1] 1.56fF
C2275 a_5743_n6391# Iref0 0.00fF
C2276 SAEN ADC13_OUT[2] 0.01fF
C2277 ADC8_OUT[1] ADC9_OUT[1] 0.01fF
C2278 WWLD[1] WWLD[3] 0.03fF
C2279 Din[3] EN 0.02fF
C2280 ADC9_OUT[0] ADC10_OUT[2] 0.00fF
C2281 VDD RWLB[0] 2.06fF
C2282 Din[4] PRE_A 0.00fF
C2283 a_5743_n6391# VDD 1.48fF
C2284 PRE_CLSA ADC11_OUT[0] 0.11fF
C2285 a_5743_n6391# ADC10_OUT[1] 0.01fF
C2286 ADC0_OUT[2] Iref2 0.01fF
C2287 ADC0_OUT[1] Iref3 0.01fF
C2288 RWL[0] WWL[2] 0.01fF
C2289 VDD RWL[4] 2.89fF
C2290 WWL[0] RWL[2] 0.01fF
C2291 RWLB[0] RWLB[1] 0.09fF
C2292 Din[15] PRE_A 0.01fF
C2293 WWLD[3] RWLB[2] 0.00fF
C2294 WWL[1] RWL[1] 22.38fF
C2295 Din[14] EN 0.00fF
C2296 PRE_CLSA ADC14_OUT[1] 0.10fF
C2297 ADC14_OUT[0] Iref0 0.03fF
C2298 ADC5_OUT[2] ADC5_OUT[3] 1.31fF
C2299 ADC10_OUT[0] ADC11_OUT[0] 0.01fF
C2300 VDD WWL[8] 0.69fF
C2301 RWL[2] RWLB[3] 0.01fF
C2302 RWLB[1] RWL[4] 0.01fF
C2303 VDD ADC14_OUT[0] 2.29fF
C2304 WWL[2] WWL[4] 0.03fF
C2305 EN ADC6_OUT[0] 0.00fF
C2306 PRE_A ADC7_OUT[0] 0.00fF
C2307 PRE_CLSA ADC5_OUT[0] 0.11fF
C2308 RWLB[2] RWL[3] 1.23fF
C2309 ADC12_OUT[0] ADC12_OUT[1] 5.51fF
C2310 VDD RWLB[11] 2.06fF
C2311 RWL[3] RWL[6] 0.00fF
C2312 RWL[4] RWL[5] 0.09fF
C2313 RWLB[4] WWL[5] 0.02fF
C2314 ADC7_OUT[0] ADC8_OUT[0] 0.01fF
C2315 RWLB[3] WWL[6] 0.00fF
C2316 WWL[4] RWLB[5] 0.01fF
C2317 WWL[3] RWLB[6] 0.00fF
C2318 ADC13_OUT[1] ADC14_OUT[1] 0.01fF
C2319 ADC11_OUT[1] Iref1 0.01fF
C2320 VDD ADC11_OUT[2] 1.53fF
C2321 RWLB[5] RWLB[7] 0.02fF
C2322 RWL[6] WWL[7] 0.01fF
C2323 WWL[6] RWL[7] 0.02fF
C2324 WWL[5] RWL[8] 0.01fF
C2325 RWL[5] WWL[8] 0.00fF
C2326 VDD RWL[15] 2.83fF
C2327 a_5632_n6430# VCLP 0.00fF
C2328 ADC10_OUT[1] ADC11_OUT[2] 0.01fF
C2329 ADC5_OUT[1] Iref1 0.01fF
C2330 ADC15_OUT[3] Iref3 0.02fF
C2331 VCLP ADC7_OUT[2] 0.74fF
C2332 ADC2_OUT[1] ADC2_OUT[2] 3.79fF
C2333 SAEN ADC6_OUT[2] 0.04fF
C2334 ADC7_OUT[0] Iref2 0.01fF
C2335 PRE_CLSA ADC7_OUT[3] 0.10fF
C2336 ADC3_OUT[0] ADC3_OUT[3] 0.03fF
C2337 WWL[8] WWL[9] 0.10fF
C2338 VDD SA_OUT[4] 1.69fF
C2339 RWL[8] RWLB[8] 0.08fF
C2340 WWL[7] WWL[10] 0.01fF
C2341 RWL[7] RWLB[9] 0.01fF
C2342 RWLB[7] RWL[9] 0.01fF
C2343 VDD ADC5_OUT[2] 1.52fF
C2344 a_5632_n6430# ADC8_OUT[1] 0.01fF
C2345 ADC7_OUT[1] ADC8_OUT[2] 0.01fF
C2346 ADC8_OUT[0] ADC9_OUT[3] 0.00fF
C2347 m1_7418_5034# VDD 0.06fF
C2348 VDD SA_OUT[15] 1.46fF
C2349 WWL[9] RWLB[11] 0.01fF
C2350 WWL[10] RWLB[10] 21.69fF
C2351 RWL[9] RWL[11] 0.02fF
C2352 RWLB[9] WWL[11] 0.02fF
C2353 a_5632_n6430# ADC13_OUT[2] 0.02fF
C2354 a_5743_n6391# ADC8_OUT[2] 0.93fF
C2355 WWL[0] Din[3] 0.00fF
C2356 WWL[11] RWL[13] 0.01fF
C2357 WWL[1] Din[0] 0.00fF
C2358 RWLB[10] RWLB[13] 0.00fF
C2359 WWL[12] RWL[12] 22.38fF
C2360 PRE_SRAM Din[8] 0.01fF
C2361 RWLB[0] Din[1] 0.01fF
C2362 RWL[11] WWL[13] 0.01fF
C2363 WWLD[1] Din[6] 0.00fF
C2364 VDD Din[9] 0.26fF
C2365 RWLB[11] RWLB[12] 0.08fF
C2366 WWLD[3] Din[4] 0.00fF
C2367 WWLD[2] Din[5] 0.00fF
C2368 RWL[0] Din[2] 0.00fF
C2369 WWLD[0] Din[7] 0.00fF
C2370 m1_4543_5034# Din[8] 0.00fF
C2371 ADC9_OUT[2] Iref3 0.01fF
C2372 Iref2 ADC9_OUT[3] 0.00fF
C2373 ADC0_OUT[0] ADC0_OUT[1] 5.31fF
C2374 ADC1_OUT[0] Iref0 0.03fF
C2375 ADC2_OUT[0] SAEN 0.07fF
C2376 PRE_CLSA ADC1_OUT[1] 0.10fF
C2377 ADC3_OUT[0] VCLP 0.88fF
C2378 RWLB[2] Din[6] 0.01fF
C2379 WWL[4] Din[2] 0.00fF
C2380 RWL[4] Din[1] 0.01fF
C2381 RWLB[13] RWL[14] 1.23fF
C2382 RWL[13] RWLB[14] 0.01fF
C2383 WWL[3] Din[5] 0.00fF
C2384 RWLB[12] RWL[15] 0.01fF
C2385 RWL[12] RWLB[15] 0.00fF
C2386 WWL[13] WWL[15] 0.03fF
C2387 WWL[1] Din[11] 0.00fF
C2388 RWLB[1] Din[9] 0.01fF
C2389 WWL[0] Din[14] 0.00fF
C2390 WWLD[3] Din[15] 0.00fF
C2391 VDD ADC1_OUT[0] 2.26fF
C2392 RWLB[0] Din[12] 0.01fF
C2393 WWL[2] Din[8] 0.00fF
C2394 RWLB[3] Din[3] 0.01fF
C2395 RWL[3] Din[4] 0.00fF
C2396 RWLB[4] Din[0] 0.00fF
C2397 RWL[1] Din[10] 0.00fF
C2398 RWL[2] Din[7] 0.00fF
C2399 RWL[0] Din[13] 0.00fF
C2400 ADC9_OUT[3] ADC10_OUT[3] 0.02fF
C2401 ADC5_OUT[0] ADC6_OUT[1] 0.00fF
C2402 VCLP ADC11_OUT[3] 1.02fF
C2403 RWLB[15] WWLD[4] 0.95fF
C2404 WWL[4] Din[13] 0.00fF
C2405 RWLB[3] Din[14] 0.01fF
C2406 RWLB[4] Din[11] 0.01fF
C2407 WWL[14] SA_OUT[0] 0.00fF
C2408 RWL[8] Din[0] 0.00fF
C2409 WWL[6] Din[7] 0.00fF
C2410 WWL[15] WWLD[6] 0.00fF
C2411 RWL[4] Din[12] 0.00fF
C2412 RWL[5] Din[9] 0.00fF
C2413 RWL[6] Din[6] 0.00fF
C2414 ADC13_OUT[0] ADC14_OUT[3] 0.00fF
C2415 RWL[3] Din[15] 0.00fF
C2416 ADC11_OUT[0] Iref3 0.01fF
C2417 WWL[5] Din[10] 0.00fF
C2418 RWLB[7] Din[2] 0.01fF
C2419 RWL[7] Din[3] 0.00fF
C2420 WWL[8] Din[1] 0.00fF
C2421 WWL[7] Din[4] 0.00fF
C2422 RWLB[5] Din[8] 0.01fF
C2423 RWL[15] WWLD[5] 0.01fF
C2424 RWLB[6] Din[5] 0.01fF
C2425 m1_6269_5033# PRE_SRAM 0.15fF
C2426 m1_5118_5034# m1_5694_5034# 0.00fF
C2427 ADC15_OUT[1] ADC15_OUT[3] 0.01fF
C2428 ADC14_OUT[1] Iref3 0.01fF
C2429 ADC14_OUT[2] Iref2 0.02fF
C2430 RWL[7] Din[14] 0.00fF
C2431 WWLD[5] SA_OUT[4] 0.01fF
C2432 RWL[11] Din[2] 0.00fF
C2433 WWLD[6] SA_OUT[3] 0.04fF
C2434 PRE_VLSA SA_OUT[1] 0.14fF
C2435 RWLB[10] Din[4] 0.01fF
C2436 RWL[10] Din[5] 0.00fF
C2437 RWLB[9] Din[7] 0.01fF
C2438 RWL[9] Din[8] 0.00fF
C2439 RWLB[8] Din[10] 0.01fF
C2440 WWL[12] Din[0] 0.00fF
C2441 RWL[8] Din[11] 0.00fF
C2442 WWL[11] Din[3] 0.00fF
C2443 WWL[9] Din[9] 0.00fF
C2444 WWL[7] Din[15] 0.00fF
C2445 RWLB[7] Din[13] 0.01fF
C2446 WWL[10] Din[6] 0.00fF
C2447 RWLB[11] Din[1] 0.01fF
C2448 WWLD[7] SA_OUT[2] 0.06fF
C2449 WWL[8] Din[12] 0.00fF
C2450 ADC5_OUT[0] Iref3 0.01fF
C2451 ADC3_OUT[1] Iref2 0.01fF
C2452 SAEN ADC4_OUT[3] 0.02fF
C2453 VCLP ADC5_OUT[3] 1.02fF
C2454 ADC1_OUT[1] ADC1_OUT[3] 0.01fF
C2455 VDD ADC3_OUT[3] 1.58fF
C2456 ADC12_OUT[2] ADC12_OUT[3] 1.32fF
C2457 RWLB[12] Din[9] 0.01fF
C2458 WWL[11] Din[14] 0.00fF
C2459 WWLD[5] SA_OUT[15] 0.00fF
C2460 RWLB[11] Din[12] 0.01fF
C2461 SA_OUT[3] SA_OUT[8] 0.01fF
C2462 SA_OUT[5] SA_OUT[6] 3.89fF
C2463 WWL[15] Din[2] 0.00fF
C2464 RWLB[10] Din[15] 0.01fF
C2465 RWL[11] Din[13] 0.00fF
C2466 RWL[14] Din[4] 0.00fF
C2467 WWL[13] Din[8] 0.00fF
C2468 SA_OUT[2] SA_OUT[9] 0.01fF
C2469 SA_OUT[1] SA_OUT[10] 0.00fF
C2470 RWLB[15] Din[0] 0.00fF
C2471 SA_OUT[4] SA_OUT[7] 0.01fF
C2472 WWLD[7] SA_OUT[13] 0.02fF
C2473 RWL[15] Din[1] 0.01fF
C2474 RWLB[14] Din[3] 0.01fF
C2475 RWLB[13] Din[6] 0.01fF
C2476 PRE_VLSA SA_OUT[12] 0.15fF
C2477 WWL[14] Din[5] 0.00fF
C2478 WWLD[6] SA_OUT[14] 0.00fF
C2479 SA_OUT[0] SA_OUT[11] 0.00fF
C2480 WWL[12] Din[11] 0.00fF
C2481 RWL[13] Din[7] 0.00fF
C2482 RWL[12] Din[10] 0.00fF
C2483 ADC6_OUT[2] ADC7_OUT[2] 0.01fF
C2484 ADC6_OUT[1] ADC7_OUT[3] 0.00fF
C2485 SAEN ADC15_OUT[2] 0.00fF
C2486 m1_2819_5034# Din[4] 0.00fF
C2487 RWLB[15] Din[11] 0.01fF
C2488 SA_OUT[10] SA_OUT[12] 0.02fF
C2489 RWL[14] Din[15] 0.00fF
C2490 RWLB[14] Din[14] 0.01fF
C2491 SA_OUT[9] SA_OUT[13] 0.02fF
C2492 WWLD[6] Din[8] 0.00fF
C2493 WWL[15] Din[13] 0.00fF
C2494 SA_OUT[2] Din[3] 0.01fF
C2495 SA_OUT[6] WE 0.02fF
C2496 PRE_VLSA Din[6] 0.02fF
C2497 WWLD[5] Din[9] 0.00fF
C2498 SA_OUT[7] SA_OUT[15] 0.02fF
C2499 WWLD[4] Din[10] 0.00fF
C2500 SA_OUT[8] SA_OUT[14] 0.02fF
C2501 SA_OUT[0] Din[5] 0.02fF
C2502 RWL[15] Din[12] 0.00fF
C2503 WWLD[7] Din[7] 0.00fF
C2504 SA_OUT[1] Din[4] 0.01fF
C2505 PRE_CLSA ADC13_OUT[0] 0.11fF
C2506 a_5743_n6391# ADC12_OUT[1] 0.01fF
C2507 ADC7_OUT[3] Iref3 0.01fF
C2508 SA_OUT[8] Din[8] 0.00fF
C2509 SA_OUT[6] Din[10] 0.01fF
C2510 SA_OUT[4] Din[12] 0.01fF
C2511 SA_OUT[3] Din[13] 0.01fF
C2512 WE Din[0] 0.01fF
C2513 SA_OUT[5] Din[11] 0.01fF
C2514 SA_OUT[0] PRE_A 0.00fF
C2515 SA_OUT[1] Din[15] 0.01fF
C2516 SA_OUT[2] Din[14] 0.01fF
C2517 PRE_VLSA EN 0.15fF
C2518 SA_OUT[7] Din[9] 0.01fF
C2519 VCLP Iref0 0.15fF
C2520 PRE_CLSA Iref1 0.00fF
C2521 ADC11_OUT[0] ADC12_OUT[0] 0.01fF
C2522 VDD VCLP 10.39fF
C2523 m1_7418_5034# Din[12] 0.00fF
C2524 SA_OUT[10] EN 0.00fF
C2525 SA_OUT[12] Din[15] 0.01fF
C2526 SA_OUT[11] PRE_A 0.01fF
C2527 SA_OUT[13] Din[14] 0.01fF
C2528 WE Din[11] 0.01fF
C2529 ADC4_OUT[0] ADC5_OUT[2] 0.00fF
C2530 PRE_CLSA ADC10_OUT[2] 0.09fF
C2531 ADC13_OUT[0] ADC13_OUT[1] 5.50fF
C2532 SAEN ADC9_OUT[1] 0.03fF
C2533 ADC3_OUT[1] ADC4_OUT[1] 0.01fF
C2534 ADC10_OUT[0] Iref1 0.02fF
C2535 VCLP ADC10_OUT[1] 0.92fF
C2536 Iref0 ADC8_OUT[1] 0.00fF
C2537 VDD ADC8_OUT[1] 1.58fF
C2538 VDD WWL[1] 0.69fF
C2539 Din[5] PRE_A 0.00fF
C2540 ADC14_OUT[1] ADC15_OUT[1] 0.02fF
C2541 ADC13_OUT[1] Iref1 0.01fF
C2542 Din[4] EN 0.00fF
C2543 Din[10] Din[11] 0.02fF
C2544 WWLD[1] WWL[0] 0.01fF
C2545 WWLD[2] WWLD[3] 0.86fF
C2546 ADC10_OUT[0] ADC10_OUT[2] 0.03fF
C2547 VDD ADC13_OUT[2] 1.55fF
C2548 ADC0_OUT[2] ADC0_OUT[3] 1.32fF
C2549 ADC1_OUT[1] Iref3 0.01fF
C2550 ADC1_OUT[2] Iref2 0.02fF
C2551 RWL[0] RWL[2] 0.02fF
C2552 WWL[0] RWLB[2] 0.01fF
C2553 RWLB[0] WWL[2] 0.02fF
C2554 VDD RWLB[4] 2.06fF
C2555 ADC11_OUT[1] ADC12_OUT[2] 0.01fF
C2556 WWL[1] RWLB[1] 21.69fF
C2557 Din[15] EN 0.02fF
C2558 ADC5_OUT[2] ADC6_OUT[3] 0.01fF
C2559 PRE_A ADC8_OUT[0] 0.00fF
C2560 PRE_CLSA ADC6_OUT[0] 0.11fF
C2561 VDD RWL[8] 2.83fF
C2562 WWL[2] RWL[4] 0.02fF
C2563 RWL[2] WWL[4] 0.01fF
C2564 WWL[3] RWL[3] 22.38fF
C2565 EN ADC7_OUT[0] 0.00fF
C2566 ADC2_OUT[0] ADC3_OUT[0] 0.01fF
C2567 RWLB[1] RWLB[4] 0.00fF
C2568 RWLB[2] RWLB[3] 0.09fF
C2569 m1_8567_5034# VDD 0.06fF
C2570 a_5632_n6430# ADC15_OUT[2] 0.02fF
C2571 RWLB[3] RWL[6] 0.01fF
C2572 RWL[4] RWLB[5] 0.01fF
C2573 VDD WWL[12] 0.70fF
C2574 RWLB[4] RWL[5] 1.23fF
C2575 WWL[4] WWL[6] 0.03fF
C2576 RWLB[5] WWL[8] 0.01fF
C2577 WWL[6] RWLB[7] 0.01fF
C2578 RWL[6] RWL[7] 0.09fF
C2579 VDD RWLB[15] 2.06fF
C2580 WWL[5] RWLB[8] 0.00fF
C2581 RWLB[6] WWL[7] 0.02fF
C2582 RWL[5] RWL[8] 0.00fF
C2583 a_5632_n6430# SAEN 0.03fF
C2584 ADC2_OUT[1] ADC3_OUT[2] 0.01fF
C2585 ADC6_OUT[1] Iref1 0.01fF
C2586 ADC3_OUT[0] ADC4_OUT[3] 0.00fF
C2587 VCLP ADC8_OUT[2] 0.02fF
C2588 PRE_CLSA ADC8_OUT[3] 0.10fF
C2589 SAEN ADC7_OUT[2] 0.03fF
C2590 ADC8_OUT[0] Iref2 0.01fF
C2591 VDD SA_OUT[5] 1.81fF
C2592 RWL[8] WWL[9] 0.01fF
C2593 RWLB[7] RWLB[9] 0.02fF
C2594 WWL[7] RWL[10] 0.01fF
C2595 RWL[7] WWL[10] 0.00fF
C2596 WWL[8] RWL[9] 0.02fF
C2597 VDD ADC6_OUT[2] 1.53fF
C2598 a_5632_n6430# ADC9_OUT[1] 0.01fF
C2599 ADC14_OUT[0] ADC15_OUT[3] 0.00fF
C2600 ADC15_OUT[0] ADC14_OUT[3] 0.02fF
C2601 ADC13_OUT[0] Iref3 0.01fF
C2602 VCLP ADC13_OUT[3] 1.03fF
C2603 ADC8_OUT[1] ADC8_OUT[2] 3.84fF
C2604 ADC9_OUT[0] ADC9_OUT[3] 0.03fF
C2605 m1_7418_5034# PRE_SRAM 0.14fF
C2606 RWLB[9] RWL[11] 0.01fF
C2607 RWL[10] RWLB[10] 0.08fF
C2608 VDD WE 0.94fF
C2609 WWL[9] WWL[12] 0.01fF
C2610 WWL[10] WWL[11] 0.10fF
C2611 RWL[9] RWLB[11] 0.01fF
C2612 m1_5694_5034# m1_6269_5033# 0.00fF
C2613 a_5743_n6391# ADC9_OUT[2] 0.93fF
C2614 Iref1 Iref3 0.01fF
C2615 WWLD[2] Din[6] 0.00fF
C2616 RWLB[0] Din[2] 0.01fF
C2617 PRE_SRAM Din[9] 0.01fF
C2618 VDD Din[10] 0.29fF
C2619 WWL[0] Din[4] 0.00fF
C2620 WWLD[3] Din[5] 0.00fF
C2621 RWL[11] RWL[13] 0.02fF
C2622 WWL[11] RWLB[13] 0.01fF
C2623 WWLD[0] Din[8] 0.00fF
C2624 RWL[1] Din[0] 0.00fF
C2625 RWL[0] Din[3] 0.00fF
C2626 WWL[1] Din[1] 0.00fF
C2627 RWLB[11] WWL[13] 0.02fF
C2628 WWL[12] RWLB[12] 21.69fF
C2629 WWLD[1] Din[7] 0.00fF
C2630 ADC4_OUT[3] ADC5_OUT[3] 0.02fF
C2631 Iref2 ADC10_OUT[3] 0.00fF
C2632 ADC13_OUT[2] ADC13_OUT[3] 1.32fF
C2633 ADC10_OUT[2] Iref3 0.01fF
C2634 ADC3_OUT[0] SAEN 0.07fF
C2635 ADC4_OUT[0] VCLP 0.90fF
C2636 PRE_CLSA ADC2_OUT[1] 0.10fF
C2637 ADC2_OUT[0] Iref0 0.03fF
C2638 ADC0_OUT[0] ADC1_OUT[1] 0.01fF
C2639 RWLB[12] RWLB[15] 0.00fF
C2640 RWL[0] Din[14] 0.00fF
C2641 RWLB[0] Din[13] 0.01fF
C2642 VDD ADC2_OUT[0] 2.26fF
C2643 RWL[3] Din[5] 0.00fF
C2644 WWL[2] Din[9] 0.00fF
C2645 WWL[14] RWL[14] 22.38fF
C2646 RWL[2] Din[8] 0.00fF
C2647 RWLB[4] Din[1] 0.01fF
C2648 WWL[5] Din[0] 0.00fF
C2649 WWL[3] Din[6] 0.00fF
C2650 RWLB[2] Din[7] 0.01fF
C2651 RWL[13] WWL[15] 0.01fF
C2652 WWL[13] RWL[15] 0.01fF
C2653 RWLB[13] RWLB[14] 0.09fF
C2654 RWLB[3] Din[4] 0.01fF
C2655 RWL[4] Din[2] 0.00fF
C2656 WWL[4] Din[3] 0.00fF
C2657 a_5743_n6391# ADC11_OUT[0] 0.02fF
C2658 WWL[1] Din[12] 0.00fF
C2659 RWLB[1] Din[10] 0.01fF
C2660 RWL[1] Din[11] 0.00fF
C2661 WWL[0] Din[15] 0.00fF
C2662 ADC6_OUT[0] ADC6_OUT[1] 5.51fF
C2663 PRE_CLSA ADC15_OUT[0] 0.09fF
C2664 a_5743_n6391# ADC14_OUT[1] 0.01fF
C2665 RWL[6] Din[7] 0.00fF
C2666 RWLB[6] Din[6] 0.01fF
C2667 WWL[4] Din[14] 0.00fF
C2668 RWLB[8] Din[0] 0.00fF
C2669 WWL[7] Din[5] 0.00fF
C2670 RWLB[7] Din[3] 0.01fF
C2671 RWL[15] WWLD[6] 0.00fF
C2672 WWL[8] Din[2] 0.00fF
C2673 RWLB[15] WWLD[5] 0.02fF
C2674 SAEN ADC11_OUT[3] 0.02fF
C2675 RWLB[5] Din[9] 0.01fF
C2676 RWLB[3] Din[15] 0.01fF
C2677 RWLB[4] Din[12] 0.01fF
C2678 RWL[7] Din[4] 0.00fF
C2679 WWL[5] Din[11] 0.00fF
C2680 WWL[6] Din[8] 0.00fF
C2681 RWL[8] Din[1] 0.00fF
C2682 RWL[4] Din[13] 0.00fF
C2683 RWL[5] Din[10] 0.00fF
C2684 m1_1095_5034# VDD 0.06fF
C2685 ADC12_OUT[0] ADC13_OUT[0] 0.01fF
C2686 RWLB[9] Din[8] 0.01fF
C2687 RWL[8] Din[12] 0.00fF
C2688 WWL[9] Din[10] 0.00fF
C2689 WWL[12] Din[1] 0.00fF
C2690 RWL[9] Din[9] 0.00fF
C2691 WWL[10] Din[7] 0.00fF
C2692 WWL[8] Din[13] 0.00fF
C2693 WWLD[7] SA_OUT[3] 0.36fF
C2694 RWLB[11] Din[2] 0.01fF
C2695 RWL[7] Din[15] 0.00fF
C2696 RWL[10] Din[6] 0.00fF
C2697 RWLB[8] Din[11] 0.01fF
C2698 WWL[11] Din[4] 0.00fF
C2699 WWLD[6] SA_OUT[4] 0.03fF
C2700 RWL[12] Din[0] 0.00fF
C2701 SA_OUT[0] SA_OUT[1] 5.34fF
C2702 RWLB[7] Din[14] 0.01fF
C2703 WWLD[5] SA_OUT[5] 0.00fF
C2704 PRE_VLSA SA_OUT[2] 0.15fF
C2705 RWL[11] Din[3] 0.00fF
C2706 RWLB[10] Din[5] 0.01fF
C2707 ADC1_OUT[1] ADC2_OUT[3] 0.00fF
C2708 ADC4_OUT[1] Iref2 0.01fF
C2709 ADC6_OUT[0] Iref3 0.01fF
C2710 ADC1_OUT[2] ADC2_OUT[2] 0.01fF
C2711 SAEN ADC5_OUT[3] 0.02fF
C2712 VCLP ADC6_OUT[3] 1.00fF
C2713 ADC14_OUT[0] ADC14_OUT[1] 5.50fF
C2714 VDD ADC4_OUT[3] 1.58fF
C2715 PRE_CLSA ADC12_OUT[2] 0.09fF
C2716 ADC12_OUT[0] Iref1 0.02fF
C2717 VCLP ADC12_OUT[1] 0.92fF
C2718 a_5632_n6430# ADC7_OUT[2] 0.01fF
C2719 WWL[15] Din[3] 0.00fF
C2720 WWLD[7] SA_OUT[14] 0.02fF
C2721 WWL[14] Din[6] 0.00fF
C2722 RWL[12] Din[11] 0.00fF
C2723 WWL[13] Din[9] 0.00fF
C2724 SA_OUT[3] SA_OUT[9] 0.01fF
C2725 SA_OUT[2] SA_OUT[10] 0.01fF
C2726 RWLB[15] Din[1] 0.01fF
C2727 SA_OUT[0] SA_OUT[12] 0.00fF
C2728 RWLB[13] Din[7] 0.01fF
C2729 RWL[15] Din[2] 0.00fF
C2730 WWL[12] Din[12] 0.00fF
C2731 RWL[11] Din[14] 0.00fF
C2732 WWLD[4] Din[0] 0.00fF
C2733 SA_OUT[5] SA_OUT[7] 0.01fF
C2734 RWLB[12] Din[10] 0.01fF
C2735 WWL[11] Din[15] 0.00fF
C2736 RWL[13] Din[8] 0.00fF
C2737 SA_OUT[4] SA_OUT[8] 0.01fF
C2738 WWLD[6] SA_OUT[15] 0.00fF
C2739 RWLB[11] Din[13] 0.01fF
C2740 SA_OUT[1] SA_OUT[11] 0.00fF
C2741 PRE_VLSA SA_OUT[13] 0.13fF
C2742 RWLB[14] Din[4] 0.01fF
C2743 RWL[14] Din[5] 0.00fF
C2744 ADC7_OUT[1] ADC7_OUT[3] 0.01fF
C2745 ADC15_OUT[1] Iref1 0.02fF
C2746 Iref0 ADC15_OUT[2] 0.96fF
C2747 ADC11_OUT[0] ADC11_OUT[2] 0.03fF
C2748 m1_2819_5034# Din[5] 0.00fF
C2749 WWLD[6] Din[9] 0.00fF
C2750 SA_OUT[3] Din[3] 0.00fF
C2751 SA_OUT[11] SA_OUT[12] 3.25fF
C2752 VDD ADC15_OUT[2] 1.53fF
C2753 RWL[15] Din[13] 0.00fF
C2754 SA_OUT[8] SA_OUT[15] 0.02fF
C2755 WWL[15] Din[14] 0.00fF
C2756 SA_OUT[1] Din[5] 0.01fF
C2757 RWLB[15] Din[12] 0.01fF
C2758 WWLD[7] Din[8] 0.00fF
C2759 SA_OUT[2] Din[4] 0.01fF
C2760 RWLB[14] Din[15] 0.01fF
C2761 SA_OUT[9] SA_OUT[14] 0.02fF
C2762 SA_OUT[7] WE 0.02fF
C2763 WWLD[4] Din[11] 0.00fF
C2764 SA_OUT[0] Din[6] 0.02fF
C2765 PRE_VLSA Din[7] 0.02fF
C2766 SA_OUT[10] SA_OUT[13] 0.02fF
C2767 WWLD[5] Din[10] 0.00fF
C2768 ADC12_OUT[1] ADC13_OUT[2] 0.01fF
C2769 SA_OUT[5] Din[12] 0.01fF
C2770 WE Din[1] 0.01fF
C2771 SA_OUT[6] Din[11] 0.01fF
C2772 SA_OUT[0] EN 0.00fF
C2773 SA_OUT[2] Din[15] 0.01fF
C2774 SA_OUT[7] Din[10] 0.01fF
C2775 SA_OUT[3] Din[14] 0.01fF
C2776 SA_OUT[1] PRE_A 0.00fF
C2777 SA_OUT[4] Din[13] 0.01fF
C2778 SA_OUT[8] Din[9] 0.01fF
C2779 ADC8_OUT[3] Iref3 0.01fF
C2780 ADC0_OUT[0] Iref1 0.02fF
C2781 PRE_CLSA ADC0_OUT[2] 0.10fF
C2782 SAEN Iref0 0.16fF
C2783 VCLP ADC0_OUT[1] 0.93fF
C2784 VDD SAEN 6.70fF
C2785 m1_7418_5034# Din[13] 0.00fF
C2786 SA_OUT[14] Din[14] 0.01fF
C2787 SA_OUT[13] Din[15] 0.01fF
C2788 SAEN ADC10_OUT[1] 0.03fF
C2789 ADC5_OUT[0] ADC5_OUT[2] 0.03fF
C2790 SA_OUT[11] EN 0.00fF
C2791 WE Din[12] 0.01fF
C2792 Din[5] Din[6] 0.02fF
C2793 SA_OUT[12] PRE_A 0.00fF
C2794 Iref0 ADC9_OUT[1] 0.00fF
C2795 VDD ADC9_OUT[1] 1.57fF
C2796 Din[5] EN 0.02fF
C2797 WWLD[2] WWL[0] 0.03fF
C2798 WWLD[1] RWL[0] 0.00fF
C2799 VDD RWL[1] 2.83fF
C2800 Din[6] PRE_A 0.00fF
C2801 ADC9_OUT[1] ADC10_OUT[1] 0.01fF
C2802 ADC2_OUT[2] Iref2 0.02fF
C2803 ADC0_OUT[2] ADC1_OUT[3] 0.01fF
C2804 ADC2_OUT[1] Iref3 0.01fF
C2805 PRE_A EN 18.07fF
C2806 RWLB[0] RWL[2] 0.01fF
C2807 VDD WWL[5] 0.69fF
C2808 RWL[1] RWLB[1] 0.08fF
C2809 WWL[0] WWL[3] 0.01fF
C2810 RWL[0] RWLB[2] 0.01fF
C2811 WWL[1] WWL[2] 0.10fF
C2812 m1_1095_5034# Din[1] 0.00fF
C2813 ADC6_OUT[2] ADC6_OUT[3] 1.32fF
C2814 WWL[3] RWLB[3] 21.69fF
C2815 VDD RWLB[8] 2.06fF
C2816 WWL[2] RWLB[4] 0.01fF
C2817 EN ADC8_OUT[0] 0.00fF
C2818 PRE_A ADC9_OUT[0] 0.00fF
C2819 PRE_CLSA ADC7_OUT[0] 0.11fF
C2820 RWLB[2] WWL[4] 0.02fF
C2821 RWL[2] RWL[4] 0.02fF
C2822 VCLP ADC15_OUT[3] 0.76fF
C2823 ADC15_OUT[0] Iref3 0.01fF
C2824 m1_8567_5034# PRE_SRAM 0.14fF
C2825 m1_6269_5033# m1_6843_5034# 0.00fF
C2826 WWL[5] RWL[5] 22.38fF
C2827 RWL[4] WWL[6] 0.01fF
C2828 WWL[4] RWL[6] 0.01fF
C2829 ADC8_OUT[0] ADC9_OUT[0] 0.01fF
C2830 VDD RWL[12] 2.90fF
C2831 RWLB[4] RWLB[5] 0.09fF
C2832 RWLB[3] RWLB[6] 0.00fF
C2833 m1_5694_5034# Din[9] 0.00fF
C2834 ADC14_OUT[2] ADC14_OUT[3] 1.31fF
C2835 ADC12_OUT[2] Iref3 0.01fF
C2836 Iref2 ADC12_OUT[3] 0.00fF
C2837 RWL[5] RWLB[8] 0.00fF
C2838 RWLB[5] RWL[8] 0.01fF
C2839 VDD WWLD[4] 0.70fF
C2840 RWLB[6] RWL[7] 1.23fF
C2841 RWL[6] RWLB[7] 0.01fF
C2842 WWL[6] WWL[8] 0.03fF
.ends


** sch_path: /usr/mpw7/Deepak/Schematic_integration/10T_SRAM_bitcell_16x1_array.sch
**.subckt 10T_SRAM_bitcell_16x1_array
*+ WWL[0],WWL[1],WWL[2],WWL[3],WWL[4],WWL[5],WWL[6],WWL[7],WWL[8],WWL[9],WWL[10],WWL[11],WWL[12],WWL[13],WWL[14],WWL[15]
*+ RWL[0],RWL[1],RWL[2],RWL[3],RWL[4],RWL[5],RWL[6],RWL[7],RWL[8],RWL[9],RWL[10],RWL[11],RWL[12],RWL[13],RWL[14],RWL[15]
*+ RWLB[0],RWLB[1],RWLB[2],RWLB[3],RWLB[4],RWLB[5],RWLB[6],RWLB[7],RWLB[8],RWLB[9],RWLB[10],RWLB[11],RWLB[12],RWLB[13],RWLB[14],RWLB[15] BL BLB VDD VSS RBL RBLB
*.ipin
*+ WWL[0],WWL[1],WWL[2],WWL[3],WWL[4],WWL[5],WWL[6],WWL[7],WWL[8],WWL[9],WWL[10],WWL[11],WWL[12],WWL[13],WWL[14],WWL[15]
*.ipin
*+ RWL[0],RWL[1],RWL[2],RWL[3],RWL[4],RWL[5],RWL[6],RWL[7],RWL[8],RWL[9],RWL[10],RWL[11],RWL[12],RWL[13],RWL[14],RWL[15]
*.ipin
*+ RWLB[0],RWLB[1],RWLB[2],RWLB[3],RWLB[4],RWLB[5],RWLB[6],RWLB[7],RWLB[8],RWLB[9],RWLB[10],RWLB[11],RWLB[12],RWLB[13],RWLB[14],RWLB[15]
*.iopin BL
*.iopin BLB
*.iopin VDD
*.iopin VSS
*.iopin RBL
*.iopin RBLB
x1 WWL[0] BL BLB VDD VSS RWL[0] RWLB[0] RBL RBLB 10T_SRAM_bitcell
x2 WWL[1] BL BLB VDD VSS RWL[1] RWLB[1] RBL RBLB 10T_SRAM_bitcell
x3 WWL[2] BL BLB VDD VSS RWL[2] RWLB[2] RBL RBLB 10T_SRAM_bitcell
x4 WWL[3] BL BLB VDD VSS RWL[3] RWLB[3] RBL RBLB 10T_SRAM_bitcell
x5 WWL[4] BL BLB VDD VSS RWL[4] RWLB[4] RBL RBLB 10T_SRAM_bitcell
x6 WWL[5] BL BLB VDD VSS RWL[5] RWLB[5] RBL RBLB 10T_SRAM_bitcell
x7 WWL[6] BL BLB VDD VSS RWL[6] RWLB[6] RBL RBLB 10T_SRAM_bitcell
x8 WWL[7] BL BLB VDD VSS RWL[7] RWLB[7] RBL RBLB 10T_SRAM_bitcell
x9 WWL[8] BL BLB VDD VSS RWL[8] RWLB[8] RBL RBLB 10T_SRAM_bitcell
x10 WWL[9] BL BLB VDD VSS RWL[9] RWLB[9] RBL RBLB 10T_SRAM_bitcell
x11 WWL[10] BL BLB VDD VSS RWL[10] RWLB[10] RBL RBLB 10T_SRAM_bitcell
x12 WWL[11] BL BLB VDD VSS RWL[11] RWLB[11] RBL RBLB 10T_SRAM_bitcell
x13 WWL[12] BL BLB VDD VSS RWL[12] RWLB[12] RBL RBLB 10T_SRAM_bitcell
x14 WWL[13] BL BLB VDD VSS RWL[13] RWLB[13] RBL RBLB 10T_SRAM_bitcell
x15 WWL[14] BL BLB VDD VSS RWL[14] RWLB[14] RBL RBLB 10T_SRAM_bitcell
x16 WWL[15] BL BLB VDD VSS RWL[15] RWLB[15] RBL RBLB 10T_SRAM_bitcell
**.ends

* expanding   symbol:  10T_SRAM_bitcell.sym # of pins=9
** sym_path: /usr/mpw7/Deepak/Schematic_integration/10T_SRAM_bitcell.sym
** sch_path: /usr/mpw7/Deepak/Schematic_integration/10T_SRAM_bitcell.sch
.subckt 10T_SRAM_bitcell  WWL BL BLB VDD VSS RWL RWLB RBL RBLB
*.iopin BL
*.iopin BLB
*.iopin VDD
*.iopin VSS
*.iopin RBL
*.iopin RBLB
*.ipin WWL
*.ipin RWL
*.ipin RWLB
XM1 net1 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.64 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.64 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net1 WWL BLB VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 WWL BL VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 VSS net2 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 RBL RWL net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 VSS net1 net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 RBLB RWLB net4 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
